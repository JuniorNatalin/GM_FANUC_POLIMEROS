��  	*��A��*SYST�EM*��V8.3�382 5/9�/2018 A��  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��  ���ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d��APPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$�VERSI3 ��� COUPLE�D� $!PP=_� CES0s!_81s! PL1> �!� � $S�OFT�T_ID�k2TOTAL_E�Qs $�0�0NO��2U SPI_IN�DE]�5Xk2SC_REEN_(4_27SIGE0_?q;��0PK_FI� 	$THKYGoPANE�4 � �DUMMY1d�DDd!OE4LA����AR�!R�	 � $TIT�!$I��N �Dd�DPd �Dc@�D5�F6�FU7�F8�F9�G0�G��GJA�E�GbA�E�G1B�G1�G �F�G2�B���ASBN_�CF>"
 8F CNV_J� ; �"�!�_CMNT�$�FLAGS]�C�HEC�8 � EL�LSETUP �� $HO30I�O�0� %�SMA�CRO�RREPR�X� D+�0��R{��Ti@UTOBAC{KU�;�DEVIC�CTI*0�� �0�#�`�B�S$INTER�VALO#ISP_�UNI�O`_DOx>f7uiFR_F�0AIN�1���1c�C_WAkda�j�OFF_O0N�DEL�hL� ?aA�a�1b?9a�`C?���P�1E�$bE�X_CN}! �� �'$� _�y �0Ya^aXsOP�TC1}bXI�PEeE�xs� TOds�RE�cuvnx�R��yp_RDY_OUj�}IA-uGW.? l 8 [p�0tt[p&U��1�3 B�� ��"; o 0�� uR�"SCA�NM� 	`-uPO�qA DF AVAILua�|��p���r������f�,� \�p�A!RD�INGByq�COEMR0T�pA�3S䇷PIR��AE A�DYs"MO� �cE' D [M�c�\�B�REV�B�~W� |�AXI� ~5�R  � �OD�Pz�$KNO^PM�;�*p���/"��� �������pX�0D`S� p E RD�_yp{ ( FSS�Bn&$CHKBD7_SE^eAG�q�"$SLOT_�H�2!�� V�d�%��3��a_ED|{p� � �"���PS�`(4%$�EP�1�1$OP��0�2�a��_OKv�UST1P_C� ���dx�U �PLACEI4!�Q͢�qbr��M� ,0$Dɦ���0�`h�EOWB��BC`T�rra�(tra��_MO�0 ����`���"F~�����PSWN#��3rZ`EN 1 �.��K�D lZ�3UL� � �[�q�� ǱM! R_gLIMka�DI�`PU�P�"س߳r軹2���TRQ��� �S_B-ORQ]6�U4a��G�_RM.őtP�3j�p؀���5�CTLĴ���%�LMñ/Ć�I\�]��ST'�\����a�Ň�Y#������BIGALL;OW� (K�":(2�0VARՄ@>�P�BL�0�p� ,Kva��P�4�� y p�X՗��CFٔ X� G�RP0+�MB�`NF#LI��Ӈ0U�P&�e$� SWITCH�HvN�P؂r�_�G�� �� WARNM�`#!W�qP�V�GNST� ��-0b/FLTR��T[��P�T��� $ACC�1a1���7�r��Iأo"��RT�P_S�Fg �CHG*�0I���T-��1��I_�T�<r��K�� x?ppj"�Q��HDRBAJ; C�����3��U4��5��6��7��� ��9{2T�C=O`S <F ����ߦ؈#92:�LLEUC]�"M��I�b��" ��1�!D:��0T}_}R   4F  <�Ft�=�)2��� 	��`T! |@� Bx�����P��_��TTO���E)	EX�q.�b����� 2 � ����"[0Ay}Rf�����sP���/� #D"�/�g�Q6���� 	����$��Bx�1P�⧢M.��P�# ޴�TRIG��% �d��8�P���`A�����e�5��� �g(:�^�R�&� t�FLEE2$�ANG AgpTBA O���1���!�Ӑ����0+P[`%�,���'����m �2b��X!;��"J;�_)R,�erCr,J>�w(
�,J�D!�Ҳ)������0fp��C�P_�POF7�(� @jP�ph�p��I9T�c�pNOMPx%3"�S]0� `T)w@&��L�� ��PA���b R�A]q�Î4�X�
$3TF^�:D30�sFSU�P�!��(c1)H�u/`1�:ESq����û�WA��cAb3�YNT��� DBG�DE7q*V;�P��tq��J�;�P�AXȀ���eT~���UF�� x3C
+ �� EGY�PI;�U*c0P�GM�HM�I�8@�FF�GSIMQ�STO�a$KEESPAT�����2����2��P_L6�4FIX
, �Lv�!dC_� �`R�Y�kSCI��hVPC9H�PhRADDdV�Q@qU�Q}W�Q�X;�_Pl"P_�P�f�Q�=�@�Rв�51]�3B�A*EUE��-�p`XF� nVGc}UGc�V�Xpc�Me�Ypcgg��!MC��.��@�SM_JB�b��a�S�g� ��e  X�b�/� �e�CHNS_wEMP��$G�0�w[��0;3�1_F�P;4�1TC1v~wT�1{��Ft�u �_V`
���lqi"uvJRS�~��SEGFRA=�ܱp�RSTy�LI9N���sPVF(�9�M �09D0��y��rl"���r b��!G'1` +�/��#��q p(��q�`����9�jH��aSIZ�od��C�TN��0h����qR�F�!,�ms߱s{���p��Rp�pL~��0p�CRC����;�ఀ�p�1q��1r)�MINI�1qr!/�߁�D�Զ�c�Cr��� �et���w����EVD����FÑ9�fsFVp�N� �a�ց��;��<c1�30�1V�SCA��0AQ�r�r1^�
2 ����t?��RGР�"?�Fțpl�FqDߵEqLEWZĮ S�����/�� t�
�v�3� I�[���P�Ez��R	0HANC~��$LG���A$fYPND���ARcP�N�Ѥq����Yse�M�E%Q�f��@`�RA��e�AZ$p�����5Oz�FCT��Π���F��L�Fp�`� ADI�OȆ����������������SG8w#���BMP�t��8�Tq1AES�Pœ��h �I4 � 	�I���CS�F5� $��Y�C�|�6�� 5$��SU9P���ARM֢ւ ��=pS@.A �<Q�CKP�##֝�#�O+�UO9�F+�F9�N+��N9��%��GRV_����DKI�DK4s��SUL9���,سDD�3��GA:�R���R��R���,�R���R��S�0���OOR��U�p� -�q� ��|�{�|��|�Q|�>��UTOOLw��� ������������‮�%�-؅�%Ғ�%�U  �M`"՟�]�XWu]ҵYO�ZO�NUk�VBk�WO�I�����X�`�H!
7 x؀���$AT��7�C�Z�Nqp�qIMG_�HEIGH�A��W�ID%P�qVT$pAC���9AA_p(����T�EXP#�D� ��CUPMMENU��8�TIT1$PROG_UD1%W!�q0BZ_~���9��UU �Ax�6;NO��ADE���� �ޯ3�p7���l�d�:���� ����AERRLV A ;c \�0��OR d�0_ID `�0�pU�N_O\���$SCYSTUIǱ�S EV�3�p��PXWO��A <r��Ke1�B ��T �TRL@= ��U AC�p�4��I�NDˀDJ\TLAY_R��A�"��kPL a�bWA����ESERVED��'A���"�U�MMY9R4"10FR}���@>����APR� 
 ?�DPOS_~@@�? F`-Ӆ��,�Ll)@y/�#8�A �A�/>2�PC@B��/#�4�PENE��0Ts�C�/#�(�L!RECi�@D�H�Cm  ?$L/3@$l#�B��`@;�pW��rN_D1�&�@RO�P�qT�?�r�� >@RIG<k�6PAUS�3�t�ETURN�2N�M[R_�0TUx0��^0EWM�r�QGN�AL}p�B$LASxˁ�3&qA$P��B$PѰ9�C�@�PCD��8�D�O�p�Y4E12�_6G�O_AWAYo2M�O�q!�g�0�D�CSS_CNST;CY4`E L(�0�;p[�BID-ѕB2*�J2�FN7@O\�2�iuBѐIj0 F� P $Z�RBlV��SPI�GPO X�I_BYɢSWT���tCHNDG�!G H� ��Gap$DSBLIO�V�eT�F^Y��tCLSr�aHFR8 OUTzY3FB�\��FEi1Z���S�DtC��IFRDOq%�^�MCpd�PP]b�R��H�W� ��D 
�tCELE���J T�@�0سINK_N��`bZ�����FHA�Fj��$:q A� vA��A�`K ��MD�LIb 2J 
�$�p�P��#��c2uC�k�c2u�cJ�c�t 2r �})tw�PdrE�	�BZ�tCSL�AVs�L�rINP��PV�P~ytA��M� %$���= س`V fV ֥FIM1�ro�sID2�s���vW���rNTV�糺rVE��tSKAI׳D����9�2i���J���� ��SAsFE�fw�_SVEXCLU�EN��ONL� ��Y�TpD��.bI_V0�^��PPLY R��cHIr��v˃_M8�}�@VRFY_�ɂMȣ��O����"�1��+�U�O�@΅cLS�0mR=$36R�P��S$SE�P{$zD!�P��q�㟔�s���Q N�0��TA�� d   �tC���AO�B�@Y��tq�L�F�R�B�����B��T��tC\�"P D �$ �BAY`�_cB�!IpK�_0��V���V� ��v���K�@QE�'RQG:�0��`PĐ ���SGҠ R ��`CUR�0�1��ʢ q ��1@wϨvߦ��UN� mT��Eʠ8dE�0K�'�$�;�,��H� �� I.�"S @� F	�K	$TOT�0�C=$��Z�:'4RTd�MPNI�"T�B���r��A-�ԴDAY4LOAD�D2$��3#�5R�EF��X�I�RU0(!�O���a`��_RTRQ5�V:�� =>�
ErJ�E��T���`�U�`"�:��D���A� .�5�W 0@A����c9p��;CM0�oSU�0����CA�Mp Xr�� NS\����IDL��W�h���S�V�GV_��|�`���DIAG���5�Yp .$Vv�0SE(�TACJ��Hq>�E�D� GrR��"�EtV� �SW{ѷ1K����2d9��`VIp9�OHO�2��PݐEtIRfGrB��¨Ï�2FqB� ��B����p�����F����`X�`>�z@B�RQ�DW��MSB�>�A�� ��i�EtLIFE �J�Y�D!TrN{�EҐ��$�y�E�C�W#�C(n@H�d@N�0Y� �1gFLA��#�OVn0�� �0GrSUPPIO�lQTr�_��ե��_X�^A��Z�W�nA����$XZ_Ab"HqY2i�Cn Tvw0C�qN� A�c�ICT�t�Z `�CACHEͶ��cץ���2�SUFFI��p��2$�3#b��� �DMSW��[� 8<�KEYIMAG�3TMC1�1�-|r�1  ���DN_D��A5��\� $[C�M� �[BD�Q�<!\MAC�2�PD�1�\A��Ĕ�P_OFT2��Q�	�ST��� �MSG�
��b�� 1�nArP\� M�1�3VN� �DV��PRDCNz������\|pFx1�ANLGF�[�1��P��A�A���b���7vc����PVIE���$1] �aBGL��$��s?�|�L��D��^:�1`STE�!T"&@\$���\$��\$�\ EMA�I�`�1ݱ��eQ_/FAUL��_$"�3�ݲQ�j@U'��0PΗ$LTT� 5� dƱI4� R�y�&2�@rP�&fc�'(��'I�,vЂ  )�TREђ?a< $>3e�S����IT5�BU!F���q���DN���'SUBj4�DC�t��|?2�DTSAV�5 w2?Ј򼁏��7��(�9P�4eORD��� �_j0�5ΰIOTT(�����P�M�u;D���8GAX�e��X�j0��3_G{�
���DYN_����b���� l�DU��MҺ���� I�T���P8��c� p� ,��"CC_R��IK���B��DopRp)�E�(�ADSPA2�BP�`-YIM�3"SHQ�c�C2�U�G����CM� IP��C��D "STH���SRr�T�"SHSD%1"SABSC'������V�d�V�P��T_D^fcCONV��Gfc��T��Vj0F{�Tpd0S� _A��SC$Ҁe��CMERĄ�AFBgCMPă�@ET��ڿ�dFU�DU�^0$���E�P҂CaDY�P,@�#�� �NOAUTO��e`:��dε�d��PS�e�C��e��Tp  �D�d?@��fH %*�aL�p�#%sLg F���E�Ct��Av��Av ��Av�Avb�Av!Av�8>y9>z{�@xJz1�Wz1dz1qz1~z1��z1�z1�z1�z2�z2J{Wz2dz�NwP~z"Nw�z2�z2�z�3�z3Jz3W{dz3Bqz3~za�[w�z3�zu3�z4�r �a���P 5�g � �$��MeINLfPLCWARMS%�� >t�RL���FAC��ST����Pj�1̚2���q�r��Jq ���EXE�Bh <H��(� ��� Me��@6��e��F{DR$�iTJ0VE��4A~�t��R~�REMM�FVq��O�VM�C��A��TR�OV��DT�0êM�XҬ��_��ª!�IND᠎�
�%0~�$DGjA��̠J ��j�DN�̠RIVx|`���GEAR�AKIOa�K����N� ����_�`���Zg_MCM~��F��;UR|bj ,�a�1�? ��]P?\߰z�?߱E���  H��1Y`i��k�)�PRA1�R�I�% X�5�UP�2� l � v3TD��P52?į ��M�G�R�S:+�BAC�Bm� TR w2�0/p)_$PROG��%�`p�Bq���IFI�� ��Y`*pw��P��T���FMR2f�n s��`qBt�L���x���������Q��哢_�qK�L�IMI� ���dC_�LvW�i�<�CLF���DGDY��LD���;�5��2���
@���G%o80J� �T�FS@H$p �P%�&�����~�$CEXI� >�&�1^@�`��'�3_�5_��9G�Q��q ��yb�SW�5ON��DE�BUGJs�☥GR��U@cBKUK`O�1� ~�PO�.�����k`����MSfZ�OORC�SMZ�=E�2 !T�����_E r /P|70`�TERM/�ys8�9 �ORI���3�t8�SMyODw24�uh�c w�v8�����UP"w�s -����r$D�ʽ�sȐG����EL�TO�!$USE�pNFIG����ʰ��: ]���t$UFR��$�`��! ̗ee�OT.`TA��P��@NSTa�P�AT�QTPTH	J�Q�`EJ �2����ART�0�����1�"���REL�
yASH�F���\�_SH�ORx`�cu� ��$��� v��u�OVR�]SyBSHI� ��Uz�b ��AYLOwPrA�AIXa�\�P�f�PERVIp'�P�
 �<a�Jq������RC��eASY1M�A�e��WJ�����EÆ�c�aU��a��A��!�e�P�[SDaORa�MF��h�����x�"�����  qA <�sHO�+�y �B�����TOC��|�ᰱ$OP� D`,P/sya�0��O,ա�0RE� RcyAXp��3]e� RZ��%�(���e$PW�RP�IM�%XR_�#VISv�o��UD�	�s" �z;�$H��!^i0ADDR6�H!�G^�1w1p1�`R�j@0@�{ H%�S F`�1Js�5�5ds�5�qsɑ�1���HS��`MN�|� `�`�"�Q�SO�LxS�@��E��f�A�CRO0��!ND�_CxS�bV54aR�OUP@ch"_
PIxP�!i!1=�҅CK� �IJp�I���Hdp�Iqp؏I~p�AC�IOAcAVED�G�C�Ey��3��} $��� _D������2P�RM_~B  P��HTTP_�`H��~ (�`OBJ�E^ar04$6�L�EMOS� �(}�2H�a_�T�R�SՐ�SDBGLVބR$KRL9HIOTCOU����G�p�LO�1�STEM�P�S�RԢ� ��� S�S�NdJQUER�Y_FLAEB�HQW�q�����0 �INCPUB?0IORf�QItib�4ja�4�jaqr��IA_C�HKCM�P �8#p+q���PxV�8RМ�pNTL�2�aR_t!~@�a�f A��7�R�h��_J��
s�S�QvIDzVA �p@03��9��Es0-vEs<u�`PRp�a �rB�1�b�q3�yTrH�Ӑ�t-uSRP�~���t�wOPw�t�����c����W�`��ĒO�THm�N�$W�Az�!�AF�1e�$BF����aWT�_��cr�9RIv�I]�TYAZ Dp�qa�UR��R_BIC>L�BYPASv�A��bm����R�`��v���Ӱ$Lh$�
$�F���C
 � ߃�P � 8�%���X��{rMA�TRIX�bC�*Lt� 3d�aFEL����0� dE�-�O�Kp/�~P�6�SHA���IZP�ATA��o$LNT�CH#ex����^C  �c��cP�1� 0հh� �2�V"l@
PD殐!հ�(  08c��1� �-�r̕ah�� D���v��������@N�aROB �F��^P�镇��U@�8�S�L�����bAL5I�b�&�DO?�o�a3PO�S�1�  =�-�BA��ف! cP��b����1�T X�$BI�A!3�a T��@�aK����F2�2�9җ�j��# �_HAN	� ��Рj����S�@2��=���j��*;AX�$aOA�yURCAN��Ax{rH�X@Sy���_B;P�B�!�q�����UBPR���q��O��"��EL�BOW�a
� 
���aL+���# ���ɱM���p<�3Y�SLICM0H)��#5E�r��PXP�#0��OSG2Ph�YSWAR$�"H�t!`��h���W��CH� �Nx� w�)�ESY9N��zSR_fAJ�3H_�pI�ES]a
uX�R��IDL�a&�cUN��S&Ѭ�0�����WNO�����'@O���a��R��R
p�_��LR��5���'����P�2 8n�R�w��Y��o�L@�~@v�{��බ�@ARGI��L_	N2P �A���a�g�o�d|�R���බ�1�� .���V⻅��鲟��LA@�sM��a��� P����w���  ��t��OT&���22F �������*!PgQ��2�M�W���m�PAI�� �� x�@t"RB â�!��	}d�Yt'|E�Y�s_|ꗨ��BJ��v������t5 ��REAI���便1u�咾HE7R�%a�� ���� ��ʤ���}�3�� ��^@UN!�o S�RM؃�>�XJ�J�(�ECKC<��`��0�Sr�Al�r��_T�a ��Ɣ�2��0ݑ��3���0REF5�q�2��10,�3��0ゔ�D�!�qETHO ��;1���`Õ�W���f$�BWh@(�IOL�j\0C����WT��bu���r�f�$C��X�"W�f�i�1#P��?�� '�c̃�TFB��ʃ'�WaMYD{r���s�$B6 �P)Cc�xu���c���l�7Vp�1]~�y���C$FR�`0{�`0W'  ��15�v4�u7��~�@H4��?;vW�pI}62���2�6�2uuW��"�WT2_	�FH&A� Ty�wX����v�'� <����	��Rt^�j� ��IoC3D_s��(���TPGLU�A�D���BINI�VcOX!�D�@AZ͡
u�W���8pߤΣ�3�z�1ׅz�2*W1�_P1�G@Q2E[3EX2B[nPSYnPbY'QPTn`�U��W �@�SnP�W�Q�V�Q�V�1T�2S�VEXT'RA1��b2���D$�� ���N�@qJR�\�3�PPEe@4De T-�FL㳽b��Z����y`PAųtdMEM^�tdP�oiPG��C�au��BZT��P�a-��U��
��
��CP�v ��O��@[d�I��@�� p��A{au� �x�C0^`CN�8��N�C�SIV/�:� S����qH&�qJ��g �Q�`�p��
�j Qr�`Nu� �aECf����f��U3�5�VE�RT���#*�����	�DLENF�H���V�ZS�MGQ�|�a�|��p���X2���Y��Z:rTOT��B���`�� B��a����{
��tא�sL�� 4� ��g����!�E+p�T�@DPf�t� $`���MjhERG�q��Vd<�C�|c0��Gķ�Z䩕��Eϒ�!�ߑ�!�!�bQ�GS��}��a��p��INO�9�&��>�p�N_XY�Idg�Zn�Gv���&� ��2�C����Pb��]���e�l@)�P�$ANALY5w�b'��	�]�Uu��b�I�c� �:a�Df�'�1��pv �  ���G��z� UpR3z�Аu������I^�BGD�v �� d �P��F	IO�V�-�c'�&и>���TAImsBOUFEX�� Q�߲u� |*`�}�[ME��a�Ir��SVq�SV~�CO�q�O~�PATJ�A)e�dk�� Be@�BOXu� @ Ҭ���_����ʁ ����^ ��^ �� ݱ)_��v �@�M��p0��$ACTC���U�PDi�A�8.ұD�# �!0Н�DZ�*�p:tOM��$TE�C ��aeq����sFL��	p$ON�a �v� A��h�3� �u �"�v��\�>@�@�� �VRWRT:�LN�TK*�ARCTOCOL�A`�� x�Z'��_ � ` �$ZPR1���B��TOK��џ�p�0���'����RV�E�������.�WĬ�@"���#PAP��
�$F�	p\.�SIB�B���e�"��B9 p4�"�\߬�ALCP�EQ�$�IO7LNK����`����q��K!� ��_���@��Pq���?�u�SLAVE{��b������������ k Xu�_�AS�A/� T��Lq�&��d$�p�RT@�	1�����~pH��5P)  pU�{����n6^ �>^ G�TRTP�K#����G�� � ��I�3q �� X��IPAD����_NE�!��LAG�!� 5 �#�q�����d$FOC�US��� ��I�TEM_AC�r�S l�� M�L0p$�p�NL7�F	 {GELA�!{E�F�4�$H8!�REP��  �G�ـ���bZ�n��N�����IRCA|0"b� � | �v�INCYC�A�8/!M�3-@3CL'I���G6�cDAY_��NTku��'��8�u��'SCAd �'�CLEAR�!�R��q@P����r%~5N_PERC�B �~!�@��C>C��7� �p��1_O�F�(>�3� �hG�qP� $w6Q2wLABـ�2��7U�B7H�@xuH<T���UJR*Q{�� � F��D�~c0@`W�2˦J7*P�c�$J8I7_AHI�E4G7�6@8KI�AAPHI�`Q�#ChGDSB_J7�J8��BL_KE�a����KARE�LM� ��XmR ON�WA���_VAV��r��1E�Ap�ty�Cq��rc�Vs��@CTR����B	c��L=D{�� x`p	��uNTD�!TdT�L��ORQcM�NTMO�\VT%�PD��Sn2 ROJ�VTOmsޏ���LG.T� ��э׿W��p�`V�WMR�W �VFD�XI�X�X���V��XP]�U�PMOD �VRf�PRf Rf`RfC`RgX_Rӱ���py~��t�LNAj�2����DE����иa�U��a�L�c�bDAU�eE�AD�aI�r�`GHv�t�� BOOz�� C/� IaT�s5tT +RE�p�LxSCRN��+Dpr��� @�RGI�� ��|��#U��u5�	S�1"W�t�d#�JGM�wMNCHL���FN�B�vK	�7PRG�UF�D�n�FWD�HLL�STP�V����<p�RS��HELHh�D� C�4b�Ec0��0�w��UF&��w ���wP8�G�y�CPO �g�wub�Mɇ�:�EXTUI�I7`&3+ 7a�r����s�����Ѱ���!	��iuѱipNwQP���TAV=��T�%PUDCS� �����*�O!�O-�Sf#K�r8�SD��xIGN�P�������ѯs�DEmV��LLRQ�#q��|���@�T͒�H��U�8$VISI��T  ���y�{����@-�o��P��;�1j�2�3'�
䳢�� � �)��T��Ku����1&LaO�Lt4A�STo �Rp��Ѱ�� ��$�в�C��@F9F��Ҷ 6�5� � � L��>R`S�����Y�2����hs_ � � $���������MC�b� �� CLDPo PUTRQLI�1RS�0����FL@���1���!)D�A��R��D�š���ORG�0����������3�Ѡt��3� �8P�Ļ��ķşSV_PT����	���p�x�RCLM�C���(ߘ�4v����MFRQq�� � !)HR/S_RU����!`@ ��k��`>�$���WOVER�c
tM��6P�EFI��%�W}���C��c \�0
�4D$M��j14?8P�!PS� �	�sP��i����U0ABP?(�8PSL�MISCN�5� d�aS�Rn�d��LPB�p� ���q�AXPR�@���EXCES8�R��M� {��� ���PTg��SCT� '� H=1��_n0���S ���/�l�MK�r�y�;T��v"B_^�@FLIC�BVpQUIREɃvP���O���V:\�ML:-�Mq� [�Dq�6 $R:S�����#MN.R��1��b�b�XuDCb��dINAUTyq�d�P@��p�N`RRa߃[�@�aPSTL�1� �4�@LOCV�RI�&0V�EX�ANG\V�����R`A�Ջ����2�0��MFRe<�|�,�6Ÿb�`��SUP2� �$��FX��IG}GHq � ��� -�Ra�$-�ӆ,��@[� �����������=�`k1ܧ@1�"P �HvڠIN��� t*MD'!�2)5&\�@$Ī�='HA@$DI<�!@$ANSW�q@$� �p�@%D	s)
�p�3n��0� ^��CU�PV~ �����l�6 LOp�0Ԙ\��$���&�2���"�&�# P�M�RR2�5�� ��!�aAu� d�$CALI��SeGt�,72�RIN��/4<$R:0SW0���j3*�ABC;D_J2SE���4!�_J3�6
�21S�P�@=���P�4�=3P�=�!CP���5J*�h�57�m�O��IM*���CSKP��$D�`$DS$DJ����Q$LUEp;EUEKG _AZtҌ�1�AEL���2��O�CMP����`R1T�a�C�%1��@�%Fv�1��H���JZ�D�SMG�� ���I'NTE����׸"U��r��Q��_�� ��$U?R�����4;Uw��IYDI�A[Q���DH?�>Pkڎ��$V90�v�$��$�@ ����$Y�1����H �$BEL��@��C.�ACCE�L\��X*��PIR�C_R��`NT<�ဳ$PS?���L  �P)f��Pgx�a�fPATH�Y�bgcbg31b�B�_���R�`�a���Q_MG��DD�a`xr$FWx� �S�e�c�R�hDE�kPP�ABN9gROTSPEE�b� S�KA��DEF���Q1`�$USE_80��P$�C���Yp�Ps�- ��YN��A<@�v�@W!�qMOU�aN�G뢰`OLRc�tINC�$�b�d��w<A�ENCS80�`��)a�R�&`IN���I1b� ��K@VEx�p032�23_U&A��D�LOWLP� �� S��ud�D���� ��P1��u��C/P+�gMOS}���MO����s�PERCH  ��0�h�̀ĆV�΃ �g�����G�Bjup`$d�CA1b#�LڔC���G,��g�b�}�T3RKׄN�AY�#� ��1b����	�F���r��MOM�r�� н ���c,7��dc��0DU@�bS_�BCKLSH_C 1b$��p��1��s��C���rM��qMECLAL�۠*�\�ӐT��CH�KS�e�S�pRTY���"�ޥ��!_�����_UM��ϩC�ܣ�aSCL���LMT�0_LРC�g!�E�)���e $�h�08��q.�j��PCԁ�H3� �e2ҥC��7�XT�P�gCN_G2N��ɶ*�SF�Q��Vjr"����Q��1bŢ�CATٮSH��G2�d�v������%2a�)�@�`P�A٤�r_Pإ��_ (@������Sѩ��Ĭ��JGe�U��R�OG|�� �TORQU\p �5�����`����` �_W땒��A�Q?Ԁ�S>ծS>�Y�e�T�I�SF��1��2��A�`�VC�P0�����1��Q������JRK�����ֱ DBL_�SM�q=�M� _D9L�Q=�GRVE�>�0�S>�S�H_�#�e`l�COSy�@y�LN���գ�P���@��p�������Z�୆�MY������TH��9�THET=0m�NK23�Sc�l�S��CBh�CB�SC��S !��pԛ�S���h�SB�S��s�GTS-A8qC�1�G����G����$DU ��F�,2�q��$ArV�Q�$NE*DBsI�ຣ�ITW$�PW�A[���k�v�v�LPHy�b<�bS ��������b���(�
��PV�V��P��V�
V�V�V��VVV H�����B���H��H�HHH* O�O�OQ)�UO�
O�O�O�UOOO�Fb����)���$�SPB?ALANCE�4���LE��H_[�SP�Q��<2��<2��PFULC@8g2O7g2���)Z1��AUTO_<����T1T2�9�R2N���R4��4WQ̑�i0G 8b�S�TS�O��@�Q/�INSEG�R��REV�6��%�gDIF|�NY1�3G6zR1ٖ�OB)Ao��H���2
�4���'�L�CHWARrorA�B����$MEC�H��(�q�A��AX���PM��F}�R P�� 
�B��Q�RO�B��CR1bU�� �i��C�Q_��T� � x $�WEIGH�pU��$�:S��I�qb�I9FTq�`LAGrl�qSr@rBILsUcODՐ��QRST�P"QRPAo�RP��P,�!Q*P�.P
�p�R�q���  2ܔ�VVD�EBUbSLZ`�R� MMY9!e@N8u�dU�$DZaށ�$�P��J� �  �DO_`A)Q� <=P�V�0��$�qN�B�R�PN(�_h�_k��p<�RO|� ��� "�T����T*A�T$`TgICKcSw@T1,`%�c��`N���0Sc��R:��q�B�e�B�e�3`PROMP�sE~<B $IR ���q��r6�UrMAI�$��q�r/u_mP�-s6@���pR3�CO�D�SFU�p_VID�_րqu@r0G_�SUFFp� hgS�q6q�bDO�g @�e�P�g�y�u�B�uPѯt3d�P�=PH]@�_FI�Q9�O�RD�Q 0P�R3"����q,`�Q6e��4 *FAL_�NAhaIpW��eDEF_Ig�W��fs��e �R�f�T�f���e���fISK ��Ka�0�d�"�cq���T4ұd�B�RD�0���SD���O0JbLOCKE u��s�o�o�g聯r�pUM�uW��t���t�� �t�r���u���t�� �r�V���s�@&Q�u W��u���s�-��x�`�P[@ք�`�` $`Wxh�g��� c �Q�GRK  � hG $���2TbX�`TMQ���^��bf���]cER'@TG�F��P�� �Q�*P� �� $GR� S�ID��B�6�D#�\�Ip6�R�3��b���sS��a/�@��.�_�9 ^@>�R��!��$�MS�K_0��� P~=Q1_USER�1��ұ�v@����1VE�LV���v@ٲ͵�AI\?�*��MT�aC��>���  �`;@�R�W�RE(Pg`���OPWOਰ�}, `SYSBUt�J�SOPA���I�TL�UK�6@P����rŃPA���téBJ�OP�pU(�f�[A�R<�Q��IMAG&��0����IM����I�N/�����RGOVCRDDb�Ű��P������@�0�"�ծBL�\�BT�2�PMCG_ED%`�@�QNt �MD��Q�R1�R,M���SLZ0���.P�$OVSL�6S\�DEX�����? nlaFF_��VR�� �p�����p���׻��RfR xh�@pTU��� @ z����EMOypRIap~
��Ep�*��  ���8AECY���� Hx=Q�@�PATUS��
aCL ��DXb�B ��o�X����QD�B���� DAa����b�}sc���Ї��X�Ei�$����������>Ph�UPR���܁PXp����T2����p�PG��? $SUBW��E���W�+�JMPWA�IT��o�LOWʭBF�aM`q�ARC�VF=q�`�Br�RE��FA�aC_CT�RO �c��IGNR�_PL+�DBTB2�PP���ABW]p��2 �Ut`��IG���`<�1�@TNLN���RT'�NOMOT�N�`�� �ERVE`��G��A�r�SP�0 � L=P�@r�g BtUNOP2�s r�R����DLY<���0a� �P�H_PKT��~�RETRIE+�<$§� c��"p;FI�� �0P� �� 2��DB�GLV��LOGScIZ�A&��KT���U#�,D�� _T�l0�BMMh0�� BE�M;RLP��FCH�ECK I���P����� 0��aiA,0I�NX0KElP8J��R��PIP��=�$ARdr�����I�OR+�FORMAT�Q���R�D	$�UX�0��� T�PL|vp��  O��SWIx@��}`AX���]pAL_ � $qAV�B7�$CCV�D���U���J3Du(� Tx�PDCK0�߂J��CO_J3&pPH@�#�#2W��/�-�P�i0 .� � �~��PAYLOA�#�$4_1+:2+3w J3AR��J875[6F3���RTIA4u95ju96V�M�PNT�3��3�3�3�3�`B��A�D�3�6�3�6�3PUB�`R�4�5�3�5�2� 
�L#���� L$PI�D*&3@aA05L.7��.7ZCJ�pnJ^KIlCR0'1��F%�F2�Q/���
�SPEED�G i"�D��d�Fd���� ���FS�H��Y���SAMP�QgaTX�G�YS��MOV_�R �Q�P��Ͳ�T�%�Vr�80�YF0ͲR [�z4�Us ٰ��U�p �[s <S�X
k�T���Z�0hd0kPkGAMM��USk��GET�I�FI�vp3�
�$z IBR
�(I$c ��R�_��q�$��fE� �hA�n�`�fLW�mv|�i1v��f2�F y!C��C�HK��=��.I_;P ��R$9(a��U�w�3�t�6�yw# ��$�( 1��pI)�RCH_�D��[�܀��|�LE@ٱ���&�8�p�+ _MSWFL��Mk07SCR�75��T3#�z��W蠁0�Y��|� ���$$C� =S�����΁Ő�Ő À�SI�!�͆ـ��:�� VMz�K �2 ΅� 0  �5�Ձ#�/� �R� R�	u�f���ŐBπ�w�������e� ؝�t���1�9���sBS蠌� 1�� <� ~�������Ưد��� � �2�D�V�h�z��� ����¿Կ���
�� .�@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖߨߺ��� ������&�8�J�\��n���I�Q`(`LM�T逕��b�  d��IN����� 	_�������v��@���Z�΁��Lp0!V� Ή��G�LM_DG 
�����ހM�_IF 
����������������+=N, 
m�u��B�����>�NGTO�L  Z��A �  $��P�FoO U� |�`Wi{�ւ a ��҂���
/� /@/*/d/N/t/�/$����/�/�/�/? ? 2?D?V?h?z?�?�?A��P@CAT�?�΅���b �SpotTool�+ �8 
V8.33P/05#��7
10412�2�2JF0'AO9�0BN�?B7D�DE�0�<GM� Global ?4 Rev0�	A�FRA�?��1DMs�_l6O`T�IV���3���AU_TOMOD�j����P_CHGAP�ONL�Op�POU�[PD 1
�� �IPM___q_�:_CUREQ 1
�S  ��{W{\g���_q����Sӂ�ق ^	�1 W{el��SW]��s�SW}`K'fHKY�_͘�_�_to�_�Pobo�o�o�^�c�Handoling�dH�U\LR�jHT;a1�o`�o�o�o�oB}c��Dispe7nseuDI{T�2
+`L/hL;oI[m ���	�'�-�?�Q� c�u����������� ��#�)�;�M�_�q� ���������ݟ�� �%�7�I�[�m���� �����ٯ����!� 3�E�W�i�{������� �տ�����/�A� S�e�wωϛϭ���� ������+�=�O�a� s߅ߗߩ�������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����������UTO� �O�C�DO_CLEAN�_
TPNM   {_�������^DSPDR3YRW�UHI�@z@�Rdv��� ����//*/�XMAX�07���a�AC&X7�qDR�q�BPLUGG7P8DS�  R�#RC	B�x |A3/�"Ox�"$SEGFP 2`�/51x�R?d?�v?�?�?�/1LAP /B>�s�? OO$O6O HOZOlO~O�O�O�O�O>STOTALj&@V}�UUSENU/0<[ �e`!_�b�P�RGDISPMM�C2`�QC1Z!@I@$<TO-O&5�8S_STRING� 1	[
��MPS�J
N�otAtPerc�h�VIsItS�af�t�RCyc�leInteru�p�TProdu�ctionSta�tusFPChu9t�X�Q  n�Mo %o7oIo[omoo�o�o��o�o�o�o�o�X�I/O SIGN�AL�UHPFr_ITEM1%#q�� �������%� 7�I�[�m���������V3�[3[y͏� �+�=�O�a�s����� ����͟ߟ���'�p9�K�]�߃WOR0 �[����c���ïկ� ����/�A�S�e�w� ��������ѿ����'PO�[FP	-��� �P�b�tφϘϪϼ� ��������(�:�L��^�p߂ߔߦ�(�DEV0���DϾ���
�� .�@�R�d�v���� ����������*�<�>N�PALT�u� ��O������������� 	-?Qcu�������c�GRIM �[���AS ew������ �//+/=/O/a/s/�/�@R鍽!1�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�?�OO)O�/PREG y�b@�/;O�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_/}��$ARG_��D ?	���a��  �	$/v	[�$h]$g�/wEi`S�BN_CONFIOG 
k;qWg�CII_SAVE  /t�ayb`�TCELLSET�UP j%HOME_IO/}~/|%MOV_�a��o�oREP�,* �;q`UTOBA�CK�`mn�FRA:\OK �,OF�`'`���OGzx� �~ FhOM��
��8�@�st���F�n� ��������ȏOE[�� ��*�<�N�ُr��� ������̟ޟi��� &�8�J�\�矀�����දȯگ��!�  �fq_Is_\ATB�CKCTL.TM�P DATE.D�x�4�F�X�j��ZFpE�Xcb ia�E�� A�sC/z  B�{e|e���GRP 3e;�` l�{OC,<�ODaOI�Pe8�J�йCܼ������"�H���X�PO_RT ��	yr0a�����OL��e�+�E�y���WRK ߻�ߎv¦�C��yc�߂�IN�Ix��uufCsMESSAG�`#�a`�wc5�ODE_D`�`�fue��\�OVc����PAUSPOS� !�k (�7�����(O ��������:�(�^� L�n�p���������U�}P��TSK  ����z�FpRCV_�ENB�`mm��UP3DT\�!�ds r�XWZDC#�qj|�STA �asaX�ISc`UNT 2�I�c �V҈�q6������% .�(��	J�4�c �: �h Eg a� ɺJ�2F�� �%D$����g4��� ľ�yB�!�f|gG�ܺ�MET� 2��PV�I�K�I�8~aI\tOI�WgWIQ2I��ڙ>���?q�@?��?���> �5�>�)�SCRDCFG 1߹%�p��e�b�{/ �/�/�/�/�/sOJ&� c/ ?2?D?V?h?z?�/ �?~�?�?�?�?OOh*O�?�$IqGR� �g ��`C�NA�`�k	It]F_ED��1l�
 �%{-�EDT-NO0z�O__pl
`�d!-Is�O��_q���G��O~_ ���E2-� Hs  l��|�L_q�P_q[���O�__qk �X�P�_
nP_b]�_��_�C3?o�O�o�nm��"Uho�oo,hao�Z4)k�of�� "U4��o�o��C5�G$�k}~ �k� ��Z���C6��� ��7�}~̏7�~���&����C7o�ߏ���}~����J�\�򟀟�C8;�{o��_�md�ϯ �(���L��C9�w�T���	�m0����������ACRr_��� 1�����eϬ���T��`@CE!K+�3��FO���"�VJ�@G�RP 2K+�X�m�y_'�ۜN ���܅�K }��������� ��~����.�� )������ ���)C�� h�B��kPu�@�P��"@+�<5?�[>���r9ȕ���?����6�ߎߞ�� r������8�>��� d�v������������ ������2����e #�~�JP}��� ����/��& w"�V����� �//=/(/6/ �/R�/v�/BT�/ '?��]?�/�?l?�/ ?�?t?�?��?#O5O GO�?kOVO{O�O\/�O �/�O�/
_�/1_�O�? �?y_4?F?�_�_�_�_ P_b_o�_+oQoOuo �o�o,ojo�o�o�o�O �O;�o_n4� �_
o���_���o 7���.��*���^o Ǐُ�����!��E� 0�"$>���Z��~ �J�\�ޟ/���e� ����t���ѯ|��� ���+�=�O��s�^� ����d�ʿ��񿬟� П9���������<�N� ���ϴ���X�j�#��� 3�Y��}ߏߡ�4�r� �����߶��ڿC��  �v�<�� ����� �������?����6� ��2���f����������$BCK_N�O_DEL  ~���/� GE_UNUS�END(:IGA�LLOW 1����j3 � (*SYS�TEM*��	$�SERV_GRP���{ POSREGƄ$���{ NU�M�
��PMU�' ��LAYE�R��PMP�ALT�CYC1�0
	AULSU��� ��LW�BOXO{RI�CUR_}~�PMCNV��}101�T�4DLIBt��2��4,n���3/E/ W/i/{/�/�/�/�- �LAL_OUT �j	7 r�9WD_ABOR"K� 0ITR_RTN� w ��3	 0NO�NSTO� K4 �38CE_RIA_�IH K5�07�~0FCFG �< �/ �1_�PARAMGP ;1;�����O!O3O�;C�  �TN�V@{�C�V@��V@�V@�V@�V@��V@�V@�V@�  �D_�D�@�@�NDiA�M�V@�V@��V@�V@��@�0D/� D�@ �@� +D3�@=�@F�@� �DY���?�@~0H�ECKCONFI�� *?QG_P�1; ��mJ_ \_n_�_�_�_�_�_�#CHKPAUS�s1j�3 ,���7�?Z=������?@�F�>r����d����~�/�_Bo� �"FoloVo�ozo�o�o �o�o�o 
D�X�O�1�?��; COLLECT_�2�jt�4�wE�N K52�rbqND�E�s!�w�7�1234567890�w�� �N��
 H�/��)@� e��,?�Q���(o���� 򏽏Ϗ�:���)� ��M�_�q�ʟ������ �ݟ��Z�%�7�I� ��m������-�t�2"�{ �@�2�@|�s�rIO $�y_�J6h�z�����6��TRP%E�_�
�L��_MOR�3�&�< U@ $B��� Q���.�πR�@�vψ���3��'��b/?�A�A{���R�K��� TP�ry)�Ma�-�?�1�Cߍ�
�u�w�k ܮ@�6dߍ���`��PDB�p+�jԥcpmid�bg���GP%�:�/  �1௴5��ap��X�#�@���H0 O9��ߜ�g�-�@ s��t��F���h����˙�̢��g��.��� y@ ���f�v�6}{�٠ud1:������?DEF *.xP��)��c��buf.tx�� ������_L64FIX ,��(���v�;c ������ 8J)n�_�������6H_E -Q�</N/``/r/�/�/@MC��2.Q(�d�%�#���2/�-��45�2A/�C:�B:�s��C�B�$?�B���CH���C2�KC�����:s�D��7D�2VD.�D��X8D�D����H6F��iE���XF%�XF��b6F�HRF�K8�9n�=�?�ƛ21�D�٫�T�4!aP�P�ϳ��1xNBN1�@CfjV@z�@4rCD����s�E�H�D���D�@F��3E�i@F�I3i>F���E��E�@H��F�@G���͑:�  >�3�3 ;�����Gnt�1��@�A5� QȦ�f¦�A����=L��<#�޵]����O��*RSMOFST (���2)�T1�D* 2��e�2�
�A��;��B��O�G?���<��M.TESTR��0_�sR�r3l��_6C@A����$���1�A
AB`2�;@1C��b��nR��:d�
�QIj�s4�]�QT_��?PROG ���R�%.�o�T>�NUSER  �u�a�q��dKEY_TBL�  Q�a|p���	�
�� !�"#$%&'()�*+,-./�w:�;<=>?@AB�C��GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������oq���͓���������������������������������耇��������������������
�i`LCK�l�U�d�`�STAT��S_A�UTO_D��a���V-�INDT_ENB� .�?P8�f*�T2v��eSFNc�5�]��GROU��6�-��Q%2���^C��CC��A�0��2`����B���=����H��z�D�;@ �I�$.��H E�W�i�{�������ß���STOP[�m�S;XC�� 27�jb��8
SONY �XC-56�_�Q�����@�9�( �А�HRC50����<�N�7`�r�Aff~��oԯ� ¯����A�S� .�w���d�����������п�+���TRL�k`LETE�� >f�T_POPр�f��b�eT_QUIC�KME|��k�SC�RE���i�kcsc�ĳa������Rc_��Uz�M��U 18Q <�܃o3߁� �<�qߋ�N�t߭߄� ���ߺ�������(� a�8�J��n������������Cus� Menu Ed�it %cus�toyn.stm��Xz��V����� v������������� A*wN`�� �����+ a8Jp������Pounce� Data�GMPNCDTA��\�'/]/�F/�/ j/|/�/�/�/�/?�/ �/G??0?}?T?f?�? �?�?�?�?�?�?1OO���_MANUAL\��m�ZCDOb9IY��b�W)TsW�O�O?�|(�wCGRҀ:�I[ B`�$�DBCOT�RIG�W��DBG_ER�RLq`;֋�Q��OL_^_p_ �AN_UMLIM���@�d�UH`DBPXW�ORK 1<�[�;_�_�_�_oo�mD�BTB_L� =���5��B4��@TADB__AWAYS�A�GCP R=���Rpb_AL�P��lb�BY�Y�Ph�n`Pw 1>�K ,��\�'��(f�n'61i_MS�IS�{k�@�@uONTIM6V��T�bv�i�
���fMOTNE�ND�h�{RECO�RD 1D�� y�01sG�O��q �1{{b$�6�H�Z��x b�������я��� ����+���O���s��� ����D�͟<��`�� '�9�K���o�ޟ��� ��ɯۯ�\����5� ��Y�k�}�������"� ��F�����1Ϡ�U� ĿN�违ϯ�����B� ������-ߜ�Q�c�u߀�ϙ߄����>�Np� ��	���?�*�8�u���IT�p�����0�`��T���x��M� Q�c����r��������0����t�8|TO�LERENCNtB���b�`L���@C�SS_CNSTC�Y 2E([ 0�arUeUb��b ������� /ASew�����UDEVI�CE 2F([ ~*1/C/U/g/y/��/�/�/�/�/1VHNDGD G(]�Cz�kULS 2H-�/U?g?y?��?�?�?�?�/WPA?RAM I�K,'�.%URBT 2-K,8p<#/�`� CI �D¯�  �I �_p�@]FTd�9IC5WA�H`@�@�\d@�@��FrD?�GKA�PH�F  \@�@�<caqAJ�B�PGD�5D�@�I�QAK[nD�bA^A�4c�M�6T�_`_ r_�_�_�_�_o�_�_�=oo&o8o�5C�,{�D0D0N�a� 	 P9M<A��+�A��,A����A��A��U2�:�`C0QB���`4�d��<�a��|%Bwq�B��0NB��QB�?>_C�o�o��ot`��? ��?� gp� �pNv �=3CUogo�Oo}� ������H�� 1�C�U�g�y�Ə���� ��ӏ���	��-�z� Q�c���=sڟ�ן ���4��X�C�|��� i����֯������ ��B��+�=���a�s� ��������Ϳ߿�>� �'�t�K�]Ϫρϓ� ����m���:�L�7� p�[ߔ�߸ߓ����� �߻�����H��1�~� U�g�y�������� ��2�	��-�?�Q�c� ��������������. ��R=va��� �������<�� %7I[m��� �����/!/n/ E/W/�/{/�/�/�/�/ �/"?�/?X?j?��? y?�?�?�?�?�?O�? 0O9?K?xOOOaO�O �O�O�O�O�O�O,__ _b_9_K_]_�_�_�_ �_�_�_o�_�_o^o 5oGo�oO�o�o�o�o �o�o6!ZlGO uo�o������ ��	��h�?�Q��� u���������Ϗ�� �R�)�;�M�_�q��� ПK��ߟ�*��N� 9�r�]��������ß ��ǯٯ&����\�3� E�W�i�{���ڿ��ÿ ������/�Aώ� e�w��ϛϭϿ�߇� 0��T�?�Qߊ�u߮���������$DCS�S_SLAVE �L�������_4D�  ���CFoG M�+����dMC:\���L%04d.C�SV���ā�  ����A ��CH��z�����m������  �m��������<���yIE�.����2�RC_OUT� N!���] �_ a}�2�_FS�I ?� &�m�������� ����4/AS| w������ +TOas� ������/,/ '/9/K/t/o/�/�/�/ �/�/�/?�/?#?L? G?Y?k?�?�?�?�?�? �?�?�?$OO1OCOlO gOyO�O�O�O�O�O�O �O	__D_?_Q_c_�_ �_�_�_�_�_�_�_o o)o;odo_oqo�o�o �o�o�o�o�o< 7I[���� �����!�3�\� W�i�{�������Ï� ����4�/�A�S�|� w�����ğ��џ�� ��+�T�O�a�s��� �������߯��,� '�9�K�t�o������� ��ɿۿ����#�L� G�Y�kϔϏϡϳ��� ������$��1�C�l� g�yߋߴ߯������� ��	��D�?�Q�c�� ������������� �)�;�d�_�q����� ����������< 7I[���� ���!3\ Wi{����� ��/4///A/S/|/ w/�/�/�/�/�/�/? ??+?T?O?a?s?�? �?�?�?�?�?�?O,O 'O9OKOtOoO�O�O�O �O�O�O_�O_#_L_ G_Y_k_�_�_�_�_�_ �_�_�_$oo1oColo goyo�o�o�o�o�o�o �o	D?Qc� �������� �)�;�d�_�q����������ˏ����$�DCS_C_FS�O ?����-� P ��J�s�n��� ������ȟڟ���� "�K�F�X�j������� ��ۯ֯���#��0� B�k�f�x��������� ҿ������C�>�P� bϋφϘϪ������� ����(�:�c�^�p� �߫ߦ߸������� � �;�6�H�Z��~�� ������������ � 2�[�V�h�z������� ��������
3.@�R{v��C_RPI*�<��� �)��e���SL�@Z�� /	//-/V/Q/c/u/ �/�/�/�/�/�/�/? .?)?;?M?v?q?�?�? �?�?�?�?OOO%O NOIO[OmO�O�O�O�O �O�O�O�O&_!_3_E_ n_i_{_�_�_�_�_�_ �_�_ooFoAoSoeo �o�o�o�o�o�o�o�o +=fas� ���G���,� '�9�K�t�o������� ��ɏۏ����#�L� G�Y�k���������ܟ ן���$��1�C�l� g�y���������ӯ�� ��	��D�?�Q�c��� ������ԿϿ��� �)�;�d�_�qσϬ� �Ϲ���������<� 7�I�[߄�ߑߣ������4PIOC 2]OK  �r�� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O��O�O��OCNUM�  �p��������RE_CHK �Q�{��A ��,8�rf_x_�Y 	 8b_�_�_���_�_�_�_o,o 
oPobo@o�o�ovo�o �o�o�o�o: Jp�_�_��Z� ���$��H�Z�8� ~���n���Ə��֏�� ڏ�2�D�"�h�z�� ����R�ԟ�ğ
�� ��,�R�0�b���f�x� ��Я������*�<� �`�r�P��������� ޿������J�\� :πϒ�p϶��Ϧ��� ����"�4��X�j�H� �ߠߺ���������� ���B�T�2�x��h� ������������,� 
�<�b�@�r������� ��������:L *p�`���� ���$Zl J�������� /�2/D/"/T/z/X/ �/�/�/�/�/�/�/? .??R?d?B?�?�?x? �?�?��?O�?O<O O,OrO�ObO�O�O�O �O�O�O_&__J_\_ :_�_�_p_�_�_�?�_ �_o�_4oFo$ojo|o Zo�o�o�o�o�o�o �oBT2d�h �������_,� >��b�t�R������� Ώ��������&�L� *�<�����r���ʟ�� � ��$�6�؟Z�l� J�|�������د��ȯ � ���D�V�4�z��� j���¿������� .�п>�d�B�TϚϬ� ������������<� N�,�r߄�bߨߺߘ� ������ �&���\� n���������� �����4�F�$�j�|� Z��������������� 0J�Tf�� z����� >NtRd�� ����/(/BL/ ^/ /�/�/r/�/�/�/ �/ ?�/�/6?H?&?l? ~?\?�?�?�?�?�?�? O O�?DOVO8/bO�O .O|O�O�O�O�O
_�O ._@__d_v_T_�_�_ �_�_�_�_oo�_(o NohO:o�o�o8o�o�o �o�o�o&8\ nL������ ��� �F�X�ro|� ��0���ď�����؏ �0��@�f�D�v��� z���ҟ����� >�P�.�t���h����� ^�̯�Я�(��� ^�p�N�������ʿܿ �� ���6�H�&�l� ~Ϙ��ϴ�VϤ����� �� �2��V�h�Fߌ� ��|����߲���
��� .�@��P�v��b�� ��`��������*�� N�`�>�����t����� ������8( n�^������ �" FX6h �l�����/ �0/B/ /f/x/V/�/ �/��/�/�/�/?�/ *?P?.?@?�?�?v?�? �?�?�?O�?(O:OO ^OpONO�O�O�/�O�O ~O�O_$__H_Z_8_ ~_�_n_�_�_�_�_�_ �_ o2ooVohoFoxo��o�k�$DCS_�SGN R�E��`�k�e��15-APR-2�2 07:29 �  �bb��06�b19 10�:40�`	p	r� S	ON��A)usQ6N��U+uq�a����y�Ӯ�~;�
;;
�cVERSION �j�V3.5.1�4	r�s�`EFLO�GIC 1S�E��  	��w�@�y�@�~��rPROG_EN/B  �t�sp��sULSE  ��u�u�r_ACC�LIM����s�!�WRSTJ�NT��a��dE�MO�|q�q�rf�I?NIT T�z�J��pb�OPT_SL� ?	�Fx�
 ?	R575�s̀�74щ6҈7҇50��1��2҄�x �|�w��TO  ����xo��|V��DE�X�d�b	p��P�ATH A�jA�\150420�22\R02\ SѓPOIהѓҐ�_VԐ���rHCP�_CLNTID y?rv�s �x��u+��rIAG_G�RP 2Y�E (<���@E�  F?�h Fx E?�`��D��A�v�BG�  ��A�������ʯ��Cf  Cy��Y�dC��q�B�i�A��mp2m6 7�89012345�6�q��@�  �A�ffA�=�qA�  AхA��HA�G���O��K��Aǥ�A�:�	q@��G��`ApG�z���A%����`B�y	qG �u��	q
9���(�A�A��
=A�˰���A��
A�Q��A�?��C����Jr������J���N����{A����?���G��K�����A�_��?��́����'�9Ͽ�E�G�A@G�:�R�A5��/K�)_�#
ϰ�����}Ϗ��ϳ��Ͽ�Pz�A�JO���?K�9p��A3\)A,��+A&C������+�=�O߽�cϰ]�W�AW��P��J?�UCK�<�4��-��%G��ߧ߹����� ���o��N������d� ����"� �2�X����� >�����������r����CM�ڱf���~�
����=�
==�G=�U>�Ĝ]���7���8��b�}7�7����@wʏ\��p��4A�p@��AhG�� �A���<i��<�xn;=R�=�s��=x<�=��~Z��;��<'A�'���?+ƨC�  �<(�Ur 4����I���UA���	p?��� ����HB�/��/=//a/s/	?)7L?S�F�"'$�/�%���V �/G������:�6��$j��L��x3A�7����u�-�b?P<�>��?��=�?�.ED�  E�  Eh�� D�0�2�?R�SzL��L�K�T��AG�;� T!��- ��a�a�z>�B���Wr�>���?b?�:�Z��=Ax���b��7���tD��D��<<o�Z3kO|MfO�O�V7�O�B�IMIC�3�t@@��C6�O
_�O.__�R_=_v_C�DICT�_CONFIG �Z`�z�t�eg�uS�STB_F_TTS�
�y��Sip�q�ZMAU�H���rMSW_C5F�P[`�  ���z�N_��L�P 3\��y P D?�e�
f%�k�g�k��?�}~�o�o�o�x�
��o�o�o(:Ht�pXj|Hw`���Hx��
����Hxg	h"�4�F�Hj�|����������̏�[�8����Z��2�D�V�4�
v�����$� ��П⟠���*�<��N�`���������Z��
�ʯܯ�x�/a0� �2�x��ɯ�c�u�w�������̵��ڿ�����"�4� F�X�j�|ώϠϲ������������2�8D�V�̴��r߄���̸x������̸ST������pB�T�f�̴�y��8���̸EE������̸45
��.� t�R�d�v��������� ���������*<N0`r�̷p����̸���Z��*<N�i(~��߲��̸���//�Zs:/L/^/̸?��/�/�
�/�/�/̶��p??*?̸��J? \?n?�?�?�?�?�/�?8�?�?�P78O(O�:OX�e�kO}O�Y�՞O�O�O�y�O�O _O(_:_L_^_p_�_ �_�_�_�_�_�O
oo�HM�6oHoZo̸�u��o�o�_�o�o�o �o	-?Qcu ��������� �%�7�I�[������DMS���������8��̴_SP"�4� F��j�|�������ğ�֟�����rT�02�D�V�Љ��v�����̸F喙�̯ޯ�̸0�� � ���B�T����$DO�CVIEWER �]�����e	 ���fr:/GMWI�ZMAN.pdf� dUU@e<�CMSP1_IT�&�  3.p����� �� �`UU`�eP  >:�S/W Inst7all� ��o� �ϓϥϷ���X����� �#�5�G���k�}ߏ� �߳���T�f����� 1�C�U���y���� ����b���	��-�?� Q�������������� ��p�);M_�`��RC_CFG� ^ĵ�!��!�������7e��S�BL_FAULTG _�
J1 N�LTTBL 1`]
 (;A,% �����/�8/ #/\/G/Y/k/}/�/�/��/�/�/�/NGPM�SK�,�e|TD�IAG aķ�ϲj�J�UD1: 6789012345r2pIf1�*�bP ? �?�?�?�?�?
OO.O @OROdOvO�O�O�O�O 	?�Ge3 ���?_>xTRECPK?]:
k4]_�7 ��?�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�O��O_vUMP_?OPTION�]FrTR�03a<u�PMESF:tY_�TEMP� È�g3B�K�p�A�p�ztUN��15�q=6Y�N_BRK b�Ĺ>2yED_SI;ZE/2' �e�x�tTAT�s�~EMGDI�rfx�q�u�NC�1cĻ ���oc�V�!�
!�d �o��Ϗ����)� ;�M�_�q��������� ˟ݟ���%�7�Iu N�`�r����������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� Ϛ�G�Q�c� uχϡ��Ͻ������� ��)�;�M�_�q߃� �ߧ߹��������� %�?�I�[�m��ϣ� �����������!�3� E�W�i�{��������� ������7�%S ew������ �+=Oas �������/ //AK/]/o/%/� �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�? �?�?�?�?O'/9/CO UOgOyO�/�O�O�O�O �O�O	__-_?_Q_c_ u_�_�_�_�_�_�_�_ oo1O;oMo_oqo�O �o�o�o�o�o�o %7I[m�� ������)o3� E�W�i��ou�����Ï Տ�����/�A�S� e�w���������џ� ���!��=�O�a�{� ��������ͯ߯�� �'�9�K�]�o����� ����ɿۿ����+� 5�G�Y�kυ��ϡϳ� ����������1�C� U�g�yߋߝ߯����� ����q�#�-�?�Q�c� }χ���������� ��)�;�M�_�q��� ������������� %7I[u��� �����!3 EWi{���� ���///A/S/ mc/�/�/�/�/�/�/ �/??+?=?O?a?s? �?�?�?�?�?�?�?/ /'O9OKOOw/�O�O �O�O�O�O�O�O_#_ 5_G_Y_k_}_�_�_�_ �_�_�_OOo1oCo UooOyo�o�o�o�o�o �o�o	-?Qc u������� o�)�;�M�goq��� ������ˏݏ��� %�7�I�[�m������ ��ǟٟ���!�3� E�_�Q�{�������ï կ�����/�A�S� e�w���������ѿ� ����+�=�W�i�s� �ϗϩϻ�������� �'�9�K�]�o߁ߓ� �߷���������#� 5�G�a�k�}���� ����������1�C� U�g�y����������� M���	-?Y�c u������� );M_q� �������// %/7/Q[/m//�/�/ �/�/�/�/�/?!?3? E?W?i?{?�?�?�?�? �?��?OO/OI/?O eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�?�?o o'o�_SO]ooo�o�o �o�o�o�o�o�o# 5GYk}��� ��_�_���1�Ko U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�C�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿ�����!�;� -�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿�ٿ�� ����3�E�O�a�s� ������������ �'�9�K�]�o����� ������������# =�GYk}��� ����1C Ugy���)�� ��	//5?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?��?�?OO -/7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�? �_�_�_o%OoAoSo eowo�o�o�o�o�o�o �o+=Oas�����_ �$E�NETMODE �1d&e��  �P�P��p�q�Q�u�U�r�xR�ROR_PROG %�z%�VE�R�� �TABLE  ��{  �@ ��]  �  ��𧏹�(c �SEV_�NUM �r  ���q� �_�AUTO_ENB�  �u�s�_N�O�� e�{�q��  *�=��J=��=��=���+<�pV�h�z��HIS���Q�p�_ALM �1f�{ ��T=��P+{���	���-�?�Q��_OUT_PUT 2g���`��P҄_ڂ�  �{;��rΪ�p�TCP_VER �!�z!=�a�$E�XTLOG_RE�Q���� �SI�Z)��STKF��+���TOL � �QDz���{A �_BWD��p�����8�_DI��7 h&e��tx�Q���STEPſ�׿�p�OP_DO�h��qFACTOR_Y_TUN��d0��DR_GRP 19i�y
�d 	ɯ����px��������glrw��qŖ�?�J �����x������x�@��B�:<B$�V@�cچ���:B?nB�1��!�����T�?�x��c�A��^?�y݊Ҋ�������\�K��U�����i�<`��>��~��P
 H�3��#���AR�1���Β<�j��i��^�I����C`}d�C��N��B�9{����UUT��|��h����E�� �����OHcEP�]��O��#Mw��K�KA������?-�g��:�6:N���9-�ڛ��������������������� �5X�FEATURE j&e����Sp�otTool+ � T����English �Dictiona�ry}�a��4D Stan�dardH ��sAnalo�g I/O	�P�7�Lgle S�hiftFq��L uto So�ftware U�pdate  0�j���mati�c Backup~
�����ground E�diting����Cam�eraT F	]�=g CellT �/�c � nrR�ndIm������� ommon� calib U}I� ���},�sh�֌��Hco� R��G� paneU o�|�Htym �select  ț�on�2M�onitor�	 иs6 t �Path�����trol R�eliabm ��9�,rner��g��L��Data A�cquis���2��( iagn�os�Q	0~�Dis�Fau�lts�bܠ�`"pense P�lug-i9$�8���( ocume��View 
���R�( ual �Check Sa�fety: ����hance�d Mirr�I�mage �Y����(Rob Se�rv�q Uk���(T1�d$�»� �&Us F�r� 1�� xt. DIO ��fiS$ [��0�@2end� E�"L>R" ���\8/7?s  9���^1�rO F0 ��	}`�UFCTN_ Menu� v#� �W�FTPw In�0fac�5_  :�ܛG� �p Mask E�xc� g81XQ��;HT�0Pr?oxy Sv�$���7{@igh-wSpe� Ski  �6�@K J0?mmunic� �ny�d,<Aur�0�0	|�U�2�conn�2	7�t@nc� ��ru 
�2���KAREL �Cmd. L�0u��  �V^�ER�un-Ti70En=vK����@�0�+� s� S/W��0��L�ic�"�"�&,v�� PogBook�(System)�	2�R�M�ACROs,,B/�Offse�H��=�8PH gri�pp c/���8PMR��Q(��u�� Mat.�H7 l�Op6# ��c�8Pech/Stop
At��Sǋb�0�$p ;��w0Mix� Q <� �ՉV8P1�Switc� �G����Q�F!.J0�u_2Tf�Pm�%h?�2f@f{il�&��	�fzQ gbG �~ka~l i Appl�@|�� %� �e�E1 p�"
���B�d-T�0�@��APCM �fun�G����GPo4$�"�d �G x�h!(Pro!� �|7PPri��F�k ��0qR Num� �#� l�@fLs50 �Adju@@	�f�W�hwp
 f,��xtatuo&���(hw��Box�	rH9�hw�) � 9��R�DM�!ot sc�ove& �-M��pem�PJ1n4 �X���p�r�!�P�!uest ԗ�,�oJ05��Q���NPX �b�B��`S�chedule0� (S=0) c�trl  qK8�~��e�!bV	o�y_�ppLibr%
�'"��7 �%~��   �=���oPt�0ssag�e �з����*&[:���� �KQ�l|X(�'CP�red  J��/�(�/I�= ��h�C TMILI�Bh���,�p�0F�irm�iX8w0�0�2Acc� �o���Ř�TX�
����@(�elynKPi����(���� GU  ����r>� Simu�la�� @@�.SPTou`P��4��O`T� �!c&~O�v. ���G�USB port� 2iPa0� a�k�� Unexc�ept� �t Z�p� /9@9�_�VC6rKB>�� �
�̠3 آ����: ���� ��p�SP� CSUI�Qۿ` �XC�M��Web�!o%	�£`Z��!bK��t�@�$�!�0VG� ������Grid��qplay }�kQ��3�� U���0iRϢ.4
 ��? ��p-20�00iC/125�L�Z@7P2 G�raphica� �����ADV-�+��C���Z@�T�'Cb� 1_��L larm C�ause/�ed�'����L sc�ii
AmrLoad�  ���[��U�pl��}LPw���� � xit ϔr@p�g3Re��Ƒ��C�3e�re�  Ck �8�0�C�*�?��pȼ rake ���� �f ����� RT/Keyb�o:Man� ��~'QUJ��H���.
�`>H,l �{Gu: .}J�P���P�   ��}�a� ycm �B2po�ri�   �"L��DCS �`./|'CX� �)������!TE �Pl��( HD�
r@�L( RAM��m��B����xcF's�7 oq: �|# 2� �|�Q~� ��!ma� N61�!.�&�� g3V�O�utput �h�T��	�
�W��EtherNeqte��$ kV0�0<���Snif%��tc��SP���ca�@�� &���FR�A�50a� ��@;�S��0�!�& Dp��Z��	��0RS =Cupomizգ��u { �1mp��P�MK�V>�`��P=k�0��P�����/�� >?|�\�E؝��}� M���`0�!;�ib0����󑦨Q�0Util���x�}���NRT�����OOn�P��l >�.9` ]Pգ��Pb"PwA/ �|�a�?  �� ��C�36  h8Òt�܁���� ��w (�`ay��I�d� ��x�� ���@f����4�a&�`%p"q�trP5/�� �Lrc��l1�xg <����@d^30eq A��y)Ģ΁W@^�tشQ@�;�0�ROS ����e���|d��0Cli�f�;�U _ 3�� i�0N�o�ڨP@-AJ�ump�J .�����So�PF���� �# �D�PEE�D OUTPUTΆ���Ę�N�/F�ILEW� H����/2�s4�G��W@Zero Do�wn�ӛS ���� �j���T�+?64MB@"c���zԋ��"FROζ+  7PϠlb<��z� !zG����t�$� 2&d����s㤂 4��1�ැ��� t�c������tr����p�,�MAIyL��Q@pz"�,�x�ࡀ� ��!�0�.�vAAdpy���L@��4s;�Q@D� 嫰GM G4� GMP1#����{�t@ABIC`X�£�D.�`Le a�rױ�� G��>�QxI���	ؐ�$�S�z�crox�v���`HWAYy�� e��@:J � ���pS4�� nt��s���-�pU�yn�.(RSS) %�l�d��`res= 4� nd�`J�$��� ��@S� �.�T���S� �A�r tex�e��;і$Lim�¿��v�o�����]>�#(�P��,=x����� SWI�MEST f4�F�!�00}q��(����_ ����<�_�S�y>��_�S�Ц(1�_c���9�o2cA\���,oNcQpAHojc+�  do�cj�����o�c�� �o�b���~�o�c��y��o�c�����o�s
�.s-��(JsC�y�Dfs���`΂s�� _�t ���sz"�P<��s�_��sϡ ���K�y�co*�� X�$��F���^@�b����k\�~�	Q�y�x�����Z0��ήd9@ ��҃�1y2����Ѓ��R��K��&��s� �B������_��aX�z���9�{���� �_�e�t�T��n�0'��ȟ�����}9$ �"���~;�>�ϐ��8�Z� B9 �v�U)��o����go��=k�䨯��)į��y��"P*����R�`�:�XsR��V��87�Ν�
�l���D�󑺈���� ̤���ֱ���ty�ܿ��L`�W���ïү,�6�b��0�R�%`�y�L�n�P|9uh�Ί�pW�S���f��i����Ï �}<������f�����a���ӀWӜ�a�~��,���)yZ�j�.U�Md�Ά���o�Ը�9�[���W@+����T������F�>y�����*��.��(��(�t�s��D�B�W9`�q||���g��g��f�*ҳ�Αխ�N����Ǭ3WL��f���珝�s���F�@�c�o�b�� �/�~�����Hx����~ज��zą����c��l����$�|�w���,�>&g?&: v� ]��Nj��X���2@�u�Q����sW���@Kˏ���T����h3� �ԙ+O�>��B7Z}�9�Tv��_��0���z���y��p��e9�o�հU��#ψ`H�/:#&��4/V#�c�<P/r#U�l/n�s�{[��/��#x}�j��K9x�/�#ȿ��5�g}�B?"����ߞR4���L?n3J3`�������4g��_�e�����4푭'�4n�����?C�񽎜O�4���,Ot&yK�jD�"&dOΆC,
/��U�Go��6��O�C`d��2�O�C��y��OԱ8_�U�J�(_JSm�@�D_fN���T�
9Uc�I�� �_R�g0��_�T��?��5� h�_vd`9o*c\k�j��Q$Wbd�B1�\on�6}�xo�c_�x���o�c8ᨙаovDc�__�d��GU�o
sH1C�C_&t��1���<^s)��Xzsd�r'_�t�sCXS��ZQ���0�?�tRsP���s�y���e;�ߝ)3��T�2P���%�sP�7��E��¨�f�DDQo�I�?�ŚᏟe�����:��|��OV���TeP���dR�l���q�GO���yq6�ƕh� ����ⓖ��Fܟ���gC�������a%N %0�R�!-3!�L��d�@�o��Ͼ`������ƨ3,֠�����ޤ��X��د�TFz9���
4ˡX��d�E�O�N�|�T�H��rQ��
P��Ϣ��R\G���9��Oڴ��Y��%5g� 0�f�����Y�+H�JĉC 9	D�fÜ�`�����`�|Ϟ�4P�y��Ϻ�t�������ϊd�}`�/��,0�T����Ήe|@�N}Y��\߆����5k3���T��ߏ�%�k@�_�ԁ@����ߖ4�ί�MQ|9 �Nu��<�E�3�X�.����ߩU3���ߩU�s���~diq���V�`��.����eϙ�?o?�#s�Z��s�
�v���W2%�"߼[�;��������o�僸����T���eN��%5 ,K4W�yK��r�%��lΎ��ߪ�>saV�B4~RC����.t���s�[�xK?�6FPz0
�3�LB4��?��9���Lvp9���s~��9U ,����,Z�k�$y*s�/2#(���N${HH/j#���d/�d�خ��/�#Z.W[o�$���/�d|���/�#;yԏ�4Ɉf07�J4LbyA[�f4A~D9`?��3C+�Z|?2tD���e��{?5qy���4:�Os�?Ί�	�rO*CMs�$OFC�_��bD1��c�~D�K3WGxO�$Zӿ�D��3cްO�C�\9P3UU��W�O��6�(_&S �y� _BSj� Y<_�Ԃ���zT�3��'ύ�:�C?�T�#3��_nD�����E�B=�_c�@�9 o�d�IHoΤg-�48oΤ4�?�Ι���:po�c=��'�o�c�l$<�o�c�����o~��v�/tMA-���o�DĩG�:t�p3�4�t&����EgTz�lnD��G/��t�1��mj����1�  H59�0��`��q21���.� R7�82  �� ��q5�>����J614  s����ATUP  K���,��545  Y�
��,�6  ����VCAM � �]�C�LIO  ?�E�h�RIa�p����h�UIF
������6H� ,��h�MSCv0�����=��}��STYL� }i�,�28  �`�I��63  `d��`h�NRE
��*@��51��p���3�@ނS�CH����߀CD�SB�  �b��P�LG  *@���DOCV�����9�CSU  �����9�����@HORS]R�0�Uk��8�����,�01���Er�EIOޝ��UJS�54�����Q4�U�wuH'd�SETZ��Rb�D�T�S�%��,�7T��9�B�MASK  �����PR�XY�@p&P��7n��_ p�pOCm��@@� ��̀l���D��> 8Nܔ���43�J6�$�@X�ϐJ53�9v0!$ӀH����-�LCH���U �ÐO�pץL�D�0̀���2J��HG�����ΐ��S�_ �������?ېM=C��. �,<�U���J�J5��}�_0��DSW  ����k�Dԑ�%s��0�ԑ�0KÐwMPRm�8� ����ɐP�r��EN  �݁�,��ɐ{^�aX���,�2��CM����"��0�f��^Ŕ�1� 1<<�ɐ��Y���I����a�ɐ�Z�J_�>�I�D���z��S���׼p�^8�?�l;,�9ɐ�6@�FR�Da�T�R3�M]CѠ`�~{�SC�o�A�G�p93��'s���SNBA  O�G����o�K._��LCa�o�;w��HL	���U��SM��Yそې�U��>��O�SPP�#3��8D�2��� ������ېHTC�=� ���TMI��� ��Ӏ���ȅ[�TPA��7�\i��TPTX � c
/�TEL�Ѡrodu<��i�ws��J8�
P�CV��duct�,�959�s_cm�p�ɐCVLO�UEC��ct\jv��FRa�com{�{VC��LOAD\��OE�\j85\�I�P��ut.ϐ+�I�v0D ��XM�857\WEBq��pc�T=� p�ro��2U�0�CG���<�IG��H�IP;GSR�IRC��a��L�p72�m���R{761�_run�	8|���AH�I����ʀY�bk.����������7H�6�2 ��p�����ˠ>�������ɐ��
p�����d�I�\n��AB���DIFw�31�f�d��681�9.f���2̀gun�J�56ɐ�Ї���9�9v=�R5��adiGѽ78�Serv�1�, P��9�=�EC��5I�I���5ȑ_swg,�@�,�.��̀8�65�wgo��8I�����\j�9�r�I�xe��Rs67U���J76��929;�8���R�5t� ��63]�!� ��J77� P�rep�7ɐeckx��F�ɐRDERȂ
��5��9I������(��65���w�R�81�) "��6�6���J879�8;\s[�NVD��<��R7t�H�FREQJ2�g��8�`�6@��l�R6��dgps ��̀�Æ�U���.�5�Gtil\�1���7P����4��9�up��8p���>�I�948���D0@Ѱ�F��CcBS!�U�TO=�p@�*�M�L�DLP!��gdg��7D�EN�DǀJNNQ���N�Nɐ725k�53�9�t��p��uch�K�GMP�� OR��IAB��
PR�ǂ3̀ing�6��ot ��P J�� ��=H II)��1��t�6 �rh ���g���CPRu�Գ�2�5\��6���ET9Sм�SLM��U����6P�@��ـL�Gene��t� �tP��t5���t847.�PdTipPio�nP �INT�Pg J8P} NPon,�=�
P����t\wtiP0G" #P��i\P*@0( Pr��� ���t������t0��t <�)%I��U��t`�um��ts_d�&��q%���tmen�&�������c2/D-��� 1�sP@�M��tU��;6,��t8��t_st`�&P��t\�)%ess0t��t��=6EN8s����t)�c&
!"7 ����Lc&29 (.�BoxPI<�PL��F\z?�z^7��/�$wge�/�+t���PF  !<7!ދfd -�6 C O�i�@P����It� �/���thk �/TK/],T�q/�*! 8�V|Ovgbk�O�+log�?�1��&��9O ��_6XI��KV���CF Spc&m T�c&
IFd&25��L��(Sa�t``6ar�&h?�$e�rl�?Z�r�6sta�_-!��U!oC�=o  � Th�& WMe�fpe�'�I7�X ��tqpg}p��	:�04�6"WT[�_F�$si�V�?�TbV_B-s1/.x_f%w�&�D?�ida��+ectsS6�,KVsuV��-tes�&�^Et�O�,nit�|x�������nG�XO��_fV4ti_?"�P�ɢ�l�b@alN�&ks2k�I�b[�NI�pon���f���I�endǯI�rcDj�l�s�H�vw���l�h��g�ůk�vrL֟�Bc\�� L��P�0�F - � 9C~��O R � ��836�v�`F (0�Y04⩖TX��bA�dS6 #1��A\�tSV"�zd�c�6m)�2\m`̟bL�Ȱ�vc2S6��o�vrg�lgruk����UP�������p�޿ ��dzM.��en ?V�0[J{96�&61 J��8�D֠`���ol�isp�f�eV�MTCS��M��7�1
�R80 �jP6q5o�U�tco��	T���a��@S���H0���$�3l�0�0��D�M (M�&mu��vi�CFu����)ph�c�֘�  �H59} �C
� 21�MI 8�2� 5 MT�O-1� P���ATUP436� @ 545��@6|�P�VCA~��CLIO���� RI�J56�O CUIF414�_ R6dP�� MSC�op\�U�0DSTYL6{28F	R663V	GCNR=<E�5E�tioj�3F�0  SCH� � �DSB���� PL�GV�e ID�OCV��ER_ D�CSU�8R6�9��ORSR���0�80Q@�0E`!EIOn�mts�54%xLѠuj983��SET"�`t�@9�@ 7t(�MA�SK"� PGRXY2�� 7
Gv  OC�MIG_=1 wel`%�"t� "�!@4A�DTP`39&H��&daddL�CHE$�`_ Os8�37_0,MH�G�dtasP S4t�#M�,MC�,0udco�"4,4�DSW6:Dt%,O�Pt%utto MPR�LBe%8�@!�EN��@e$\vgvO160DIF/ �PCM�04 R�  0�5� "E01\h 2e$,� "�\$�5�5�0�j70�O PRS$�R5Ҥ \@@9e$704.FRD�7Int  MC�4�#�S��#H933�p� NBA�S5.�BSLC�r0P� �HLe,SMUvAc�Bu`QpPu	aP`2,�@REw4\a�HTCU�TMI��@� " �$�TPA5���Q�TX"� TEL��4a| 2�$��J�8$��6 NT[ "@ 95uE(�Q8�Pe$�SUECE$� ο UFR��#VC��E�рO�8� I�P�fl� SUI�"�g�RCSX�5�25/ WEBUi���`QTUed�ARK62u � � G�e��aIGde"D�J? IPGS&YI�RC�djd?Hs72%#R765\�a��u,C��� ���lR7% Eaq�#F� �186�m"J9TUFron< rLib,0e$x���R\awm�"veMF�0CAB��,SR53Eon\�o8E�BPwmfO26e$<c� �c{R5�erio5@r\uE�R71�we ��D75��poq5 d%��@uYП0B�ien�@2�$�� �M�f0EZ��m��q67uMN0!6�y���8$Eink��5�VI/? B%j�P80!7J5/ �R57�ux�`e$J�8>���Oh��B�X�P�� rcli�0%ECO�PR8�1%����$�po8u71bNVD$܌��U_at�BEQ���8�wr_��65̄6�%l�@�5��BbpU5�RB %ɳ���BEse�Ra7�Uh��U�R84�4cu0p%v�D]0uR H/�F��CBS�enuNO�CTOU�0F���)�V�LP�\�rs_ p�$ �@ N�N\s"�e$�vs\hQ54-���GMP$ / IA�Bed��@fin"��6�u�@? S,��	PHԥs�����M�6��H���$�C{PR��gmvz  ��F�0�D�0bET�S�dY�QLM$a�����$�cP%�3G�eneR�s\s�%�X�q�l�q�|�q�plibpɜ�q��q� ��q�̲q�ܲq����leq��>`q����<-�q�tn.p ��� p�LR��l�p��� 8p�����rop��� ����q����=aqȌ8�Q��qui��1�q�m�/ڼb��md. p�|�q�BqȜ�����qȼ��ɭ�q�ntu��ʬ2�� Q��p�k =�qȜ1��1a�m�,B<��r�g1.vp���I2��`�4����r��`������p�fy.���cN��tn��d.�AX_�
 ��NU �$M���S�p�_CO�
AR �$p�3] 6p�S;ec�  !�@��-p/�- R�
i�za��\r�mq��S4�atiڜ"A��C�
L�rc\f �#1�ϡ
�P��S�Ȩ,p����-Q��\mhpς�4/ f�_ڼ��������f�h�0!�3��W�-�?�"Q�m`��'��0�)���:pinoʬB�(LB �	�� ��$���\0@�R�d��tp����S/��x������mlan�������FOXOjO\gm�:l?~?�)2�?�?Q�J�_�_:u^�p߂�p�ߦߘj�afe0_ B_T_v/�/�/`�?�? �?�O�O.O`_r_�_B�Vw�O�O�O&�o�O��O�O�O__ mcel�������_�_ o3EW)�yo� �����Q������pg�1�C�U�g��y� mdioʜ� ���o�o�o�o ,}��Ο:����0#�5�G�Y1pr�j�� ����ҏ����/�/��zpλ�/?`�r�����t_��������ȯ`گ,}�.�0�vaN��`�r�$?6?H?��ms�*o.o�jgNo`oro��o�o�o  wiz _���������(�:�L��,n�|ߎߠ߲�����vi�������ܰ �  �STD9�LA�NG��zvis ��l���l� �1L��Q a|�4-�d��x<!gmpn ���L�XͰntr�0BT	ܱ�dv����er H]���\�x�0auto��p��
	tock&T
a.O&����8&M0ȸT�/��sy�r "8��yrs��	wtia�  !S��� .8&spk-� Sg(!&R R�NH57RI�N�&gI8d Ra�8&II)��P&p�d�'"RMTX�PLl�@ets�O&" #18&! r'd<0.fdS�imi��64�3S0 H6L66�20$F7' H7�3F06S8-J8�7t&,@8'65F3e0S5P@L673/F�9h@HHC&61�G2�-J1�F1EK27�2"G6�K�66�@�RBTi�84�OPTNf@68� DV-AETH663�DU2�@DUNT "DUSLMTDUBET�I)~W��DUmt\�s�XVFS\sl�mDUr�ET�P�V!� n1DUPosi�DUtilfPET0|�Au_ N100DUson�ETes,OV� "6 ETh�Upo�V1�XnIh! h�8�VualDUxe�sDU��ea1ETgl@PdfDrf P� `e�0DU�ET73~W܌�DV73.dfam�f- AMXfviqcdf�ePRI�V�ngcgIn{fe,� vm`�V|�Xfx\-a�VX"OVF 0DU��0�f95.fpfe<�w<2DPN ���`
�}PL�895�OP
�den�P
�a�rt+��0O��0h� "NO��	��px{`:�}�Mome���CO�APgP
�"Lyo�p
�A (C�nt A�A�s���	�t\cǆ���!� ���p
�C-f̷`
�on��<�oted >R3��upNX��pCX�le�x X�5�,X��PxX��"�x\cxX��TP�p��2�cfl��mE��Rq����Ė�ş�c�Rem���<2��a����897�@�LAS���0h{�L"I�\X�SR����r��w�  q X���thaۖ9
�X�- C��10Qe��J�%�P��d�p�X�ont.|�ed����pd�,r��%1��r�Lin�o�org�BY�k���e T�d�q��r��rq�cltȶ�19��p���19�008�dia8����uq�r�G M���p'�p"�� @7�)�\swܖG������J @ܟ" ���D�|���o�}��guif��p���Q��51�Rv@�ar-y/�J6�d'�}P�o�ally�GZ��to�@���W�TX�ϊ�sg���0{�DL�3��Կ��g�P��������Q�f�tsk���� Se��mD������
�	a�l�9�@`�|P|�J95 �n{�a`ǿ�������2j���c�ap{� �CD��o7adi��(S�E� $�|ƅ1�K�-��~P�Q���(����2��hi�s�L��l�� cd ���������wn�L��1�S012��74���l�{�D�C\И�y{ L��CD (|� H�ߢߴ߮h ��BTfkh\�� ��4���\�zd��π��- �d� 2���Prim8{��21�1F}�ss�=0O�G�����RS�sur�������pr�� � ���ɢ�v�73ngl`�nr�ang��TNtM��t'�g "��0r	�q��ad��5 c�xb��!0��D!��pfc�ir�pe�ce���Im��0�H590��a%6RS֤?�/t�wnmi��"EMg�(��r.v�� ��2<)p}��� To�0��R8J`��Ł��1 c(M������cp��BUI���Rm5mb��iMK&/�gr�'� �67b�t�FSqW@�+���7\f�ƹR����j96;�h�ٟOT\���h:f_8֐/^�_re'�(�'�ut.w�t��P/�__��O=�_en���j9@�Qocn�_�n4w旀?��P`l�i�b��
��&����!�����fx���%w�E��&�JĨ���oMb\v4�CV><?  vcfo�(��c99^���H�$FEAT_�ADD ?	������   	ux"�4�F�X� j�|�������ď֏� ����0�B�T�f�x�����DEMO �j�    ux˝��ӟ ���	�6� -�?�l�c�u�����Ư ��ϯ����2�)�;� h�_�q�����¿��˿ ����.�%�7�d�[� mχϑϾϵ������� ��*�!�3�`�W�i߃� �ߺ߱���������&� �/�\�S�e���� ���������"��+� X�O�a�{��������� ������'TK ]w������ �#PGYs }������/ //L/C/U/o/y/�/ �/�/�/�/�/?	?? H???Q?k?u?�?�?�? �?�?�?OOODO;O MOgOqO�O�O�O�O�O �O
___@_7_I_c_ m_�_�_�_�_�_�_o �_o<o3oEo_oio�o �o�o�o�o�o�o 8/A[e��� ������4�+� =�W�a�������ď�� ͏����0�'�9�S� ]�����������ɟ�� ���,�#�5�O�Y��� }�������ů���� (��1�K�U���y��� ����������$�� -�G�Q�~�uχϴϫ� �������� ��)�C� M�z�q߃߰ߧ߹��� ������%�?�I�v� m����������� ��!�;�E�r�i�{� ������������ 7Anew�� ����3 =jas���� ��/////9/f/ ]/o/�/�/�/�/�/�/ ?�/?+?5?b?Y?k? �?�?�?�?�?�?O�? O'O1O^OUOgO�O�O �O�O�O�O _�O	_#_ -_Z_Q_c_�_�_�_�_ �_�_�_�_oo)oVo Mo_o�o�o�o�o�o�o �o�o%RI[ ������� ��!�N�E�W���{� ������Ï������ �J�A�S���w����� ����������F� =�O�|�s��������� �߯���B�9�K� x�o����������ۿ ���>�5�G�t�k� }Ϫϡϳ�������� �:�1�C�p�g�yߦ� �߯���������	�6� -�?�l�c�u���� ���������2�)�;� h�_�q����������� ����.%7d[ m������� �*!3`Wi� �������&/ ///\/S/e/�/�/�/ �/�/�/�/�/"??+? X?O?a?�?�?�?�?�? �?�?�?OO'OTOKO ]O�O�O�O�O�O�O�O �O__#_P_G_Y_�_ }_�_�_�_�_�_�_o ooLoCoUo�oyo�o �o�o�o�o�o	 H?Q~u��� ������D�;� M�z�q���������ӏ ݏ
���@�7�I�v� m��������ϟٟ� ���<�3�E�r�i�{� ������˯կ���� 8�/�A�n�e�w����� ��ǿѿ�����4�+� =�j�a�sϠϗϩ��� �������0�'�9�f� ]�oߜߓߥ߿����� ����,�#�5�b�Y�k� ������������� (��1�^�U�g����� ������������$ -ZQc���� ���� )V�M_���  �����/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w�������  ����ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I�@[�m������������͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ��������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7�I[m�����$FEAT_DEMOIN  �������I�NDEX�����ILECOMP k���!��� SETUP2 l%�%"�  N� P!#_AP2B�CK 1m) � �)��/�+%z/�/� �/�/� y/?�/2?�/??h?�/ �??�?�?Q?�?u?
O O�?@O�?dOvOO�O )O�OMO�O�O�O_�O <_N_�Or__�_�_7_ �_[_�_o�_&o�_Jo �_Wo�oo�o3o�o�o io�o�o"4�oX�o |��A�e� ��0��T�f���� �����O��s��� ��>�͏b��o���'� ��K���򟁟���:� L�۟p�������5�ʯ Y��}���$���H�ׯ l�~����1�ƿؿg� ���� �2���V��zϠ	χϰ�*)^ Pb/� 2w 
SYSS?POT.SV��c�{*��TEM*�-� %-�T�>���π�ߤ߱� 8B���f�EALw߉���0�;���[�����@� ������7�p�LSCH���9�<� ��c�����(�`������h��IO������@;�!��k���0����7��*.VR u�" %* �Km�P�tPC��FGR6:���`� TX�)/� �H/U)�y/;�*c.F/�/%	���!�/�(h/�/�+STM�/2?��1P?"]9�/�?�+H?�?�C7�1�?c?�?
O�&GIF�?:OE5&AXO�?8|O�O�&JPG)O�O�E5�A�OkO __JQS/A_o��CSD_��O
JavaSc�riptm_�OCS�S�O�_E5�Q�_�M�Cascadin�g Style ?Sheets�_C��AZ*.BIN� �_a�FR5:�\4elo�IAut�oZone .bin fileo,iDAT;oMo_g�a8�oo�bdat�oc��ARGNAME.)D�ob�H0\<�o�TQlt})lpDI#SP�`uX:� ���u�q��
KVAREEG��grD�p��O��d�POSw��܏cvȏ����-�;�	GREG��`�n�hq L�
����d�u��ax�П����5�t�TPLsIN�j� %hq�T��$���d�TPEINS.XMLį�쟂�گ��%Cu�stom Too�lbar�t�PA?SSWORD��aΏFRS��]��%�Passwor�d Config<��u�WPAT�`�뿦���2� %�BU:Spot �App Proc� pa!�k�gmc1�.v=�G^d�|�}υ0�Fp��=�d�f3g*k���%�� �~+�%Wiza���"G�gmpncd�ta����lՄߪ�Pounce DJ��Z�GMWIZLO�������ߞ�|�@�L�og��D�atf�m t߆�t��v�0�A��tion GRS4��L�MP�������&�8�MHPLG?����h�����x{���� ���� ��r���=��a ����&�J�� ��9�2o� �"��X�|/ #/�G/�k/}//�/ 0/�/T/�/�/�/?�/ 0?U?�/y??�?�?>? �?b?�?	O�?-O�?QO �?JO�OO�O:O�O�O pO_�O)_;_�O__�O �_�_$_�_H_�_l_�_ o�_7o�_Homo�_�o��k�$FILE_�DGBCK 1m����`�� ( �ΐ�UMMARY.D9G�oh�MD:�o�L�Diag SummaryCONS%��o�D:X�'q��s?ole lo¿��?TPACCN���%��#uTP wAcc��tin��F��6:IPKD?MP.ZIPL�|��
d���$u4�Exc�ep�ᡏR� pME?MCHECK�u�$���Memo�ry��P�ބ=)�RIPE�������3�%k� ?PacketN᩟�]����k�ST����������� %}��StatuM�ܜ	F��p�������0��qmment� TBD��Y�ep��)ETHERNE�������4�'qEthernɐ���ur��5�ܰ��DCSVRF���������=�{� verify all���\���(v�DIF�F������;Ϻ�иd�iff=���{�CHGD12��+���� R����|�~�2�ϝϯ�D� q��k���GD3:�8!�3��� Z����~�UP)�ES.�)��FRS:\��M���Upb�e?s ListM�J{�PSRBWLD.CM|��8��O��9�PS_ROBO�WELү�� �I�r�*���N�1�L�N_et/IP��aΟ�u��rh)@�G�RAPHICS4�DJ�3�E�W�%�4D Graph�ics File�N�v�Ƿ�f�SM�q�2��V1�/�Emailw�p��{l,�NOTI���5G�3�Not�ific]� r�����SHADO�W���b5�S�hadow Ch�ang��r���~�RCMERRZ�?Q�5��CF�G Error �Det{ � ��ި�CMSGL�IB���l/7��/%H�m���m/% �t)X ZD#�/U/��/1�ZDːad��/,�l)� I�RDG_REPO�R*��/�/�/%�iR,qno2 R�eporo� ���PRCSW�c0j?Q?c?�?�2Sp�ot App p?rocess����9|�(O�?�?�-e;%Oog HO߅�0MP�?VOhO�OT��MH PlugsinOoɉ�X:E��C�O�O�O_ h%�_�O<X�VAR���z_b_t_�_�$ V�archgB�ba�se	o�TPDR�A�O�_�_�o 5Oc ��8�ox�tA�)���o�o��o5@���o72F'd�o ���M�q� ��<��`�r���� %���I��������� 8�J�ُn�����!�3� ȟW������"���F� ՟?�|����/�į֯ e����������T�/H�$FILE_8�{PRG���C����n��MDONLY 1�m��5@ 
 ��:B_VDAEX?TP.ZZZ`���近l6%NO Back f��9 ¿s����I� ؿm�6�zϣ����V� ���ό�!߰�E�W��� {�
ߟ߱�@���d��� ���/��S���w�� ��<�����r���� +�=���a������� ��J���n���9 ��]o���"��~r�VISBCK��|����*.VD���FR:\� I�ON\DATA\��5BxVision VD�@N ������q� /�</�`/r//�/ %/�/I/[/�//?&? �/J?�/n?�/?�?3? �?W?�?�?�?"O�?FO �?�?|OO�O�OmO�O eO�O�O_0_�OT_�O x_�__�_=_�_a_s_�oh�MR2_GR�P 1n����C4  B��P	� ��OoalL`E�ˀ wo�kL`OH�cEP]��O���#M�˫aKA���m?�`�ol�L`:6:N=��a9-��e�m�A�  ){BH�IcC`}dC��=NGqB�{Oul�Kdq�}L`@UUT�U~��k��Ka�>FD�>�d��>D�=��=��1��`�H�$:��=:���:.�	:sf�:�Uf�8���5�n�Y���}���l_�CFG o��T ����&���NO ���F196843 �   �RM_C�HKTYP2������P�������q�OM�w�_MIN2��S�������Xr�S�SB؃p����Mf֟�U͓����m�TP_DEF_�OW��T��#�I�RCOM|�.��$�GENOVRD_�DO����\�TH�R�� dx�da�_�ENBM� a�R�AVC+cq���� �of�}`�}�EӤ�G
��F�/lG�,Л��#��RK`������f)�gri�����OU.`w2l��P_h2�P�8��m��Y���ͿϿ/  C���	ϛ�lA��XB�1�B�pa�:�biz�� SMT�ȣxϩ>`̐��$�HOSTC؂1y����_ 	��������V�F�e:�k�}ߏ� �߯�Y��������+��,��	anonymous/�]�o����� �������%� G���6�H�Z�l��ߐ� ����������1�C�  2DVh�������� �����
.@ ��dv���� �//*/</�� ��/��/��/�/�/ ?I?8?J?\?n?�/ �?��?�?�?�?�?E/ W/i/{/}?WO�/�O�O �O�O�O?�O__0_ B_eO�?�?�_�_�_�_ �_O+O=O�_Q_>o�O boto�o�o�oUo�o�o �o'o(o_L^p ���_�_�_o�% Go$�6�H�Z�l��o�� ����Ə؏�1C � 2�D�V�h����� �ԟ���
��.�@� ��d�v����������������*�����E�NT 1z~� ?P!PLC;�����!124�.11.240.31���!��̿���� 92.168.1.54Ͽ��� ڼ8���\�n�1ϒ�U� ��y��ϝ�������4� ��X��|�?ߠ�c�u� �ߙ��߽����B�� ;�)�g��_������ �����,�>��b�%� ��I���m����������(��L	QUOICC0X4���5g���!1�2�e	��E�Fi Router�H�!���PCJOG�s���鴑0qfCAM�PRT����1��RTR8//&/��/M�NAME �!Y�!ROBO�/�/S_CFG �1yY� ��Auto-s�tarted��FTP��1���� J?�n?�?�?�?�?S� �?�?�?O3?!O�?XO jO|O�O�Oq��/
?? �O0OR?_A_S_e_w_ >O�_�_�_�_�__�_ o+o=oOoaosox��� �����_�o&_' 9Koo���� �o\���#�5�G� �o�o�o������o׏ �����1�C�U�g� y��������ӟ��� 	�P�b�t�����u��� ������ϯᯨ��� )�;�M�p�򯃿���� ��˿ݿ$�6�H�%�\� Iϐ�m�ϑϣ�j�`� �������2�3���W� i�{ߍߟ����
�� ���R�/�A�S�e�w� >ߛ��������� �+�=�O�a�s����� �ߌ�����&�' 9K�o����� �\��#5�/�� _ERR {��*EUPDUSI�Z  � ^����l>�WRD �?�%���  �guest �����//�$�SCDMNGRPw 2|�%o����� ������ � Kd$ �	P01.00� 8��   �A  %  
Vc Ϙ }���� ������������h� 1�� ����X�- � ��'�  k�����/�y�'��E���R��[��/�� � Yӝ�+ 
����/��{� �0-� �j� e� �$?؄8%���3sZ�/�/��/�/=+_GROU�O }df 1"	�G!�#�8QUPD � ��l�48@T�Y�@dWTT�P_AUTH 1�~d <!i?Pendan+'�N���0 !K?AREL:*�O�O�MKC�O�O�O�@�VISION �SET@Q_(_� �Bh_V_�_�C�_�_�_ �_o�_�_9oo"npDCTRL d�"�h
� �F�FF9E3Eo���FRS:DEFA�ULT�lFA�NUC Web ?Server�j�a VsA��Xl!3E�Wi{SWR_C�ONFIG ��S+ f�oUIA�_CHKCMB s2�S'� �d$� !ROB�O�m�Xe@@y��Xb"�g X`B�4� f"���f�e����@z2�D�V�h��c!ُ��#���Ǉ �Տ������/�A��S�e��rDEBUG ��{
�B�&���a�N�5�r��DE�L ��{��8�?�q������vELB��ǥ{�%�����Ä ˟ݟo��� ,�>�P�b�t���򿪿 ��ο�q��ϧ�:� L�^�pςϔ�%߸��� ���� �ߣ�6�H�Z� l�~ߐ�!�������� ����2�D�V�h�z� �������������
����.�@�R�d�v��wF�OBJ 2��|��*�PQ�izQ�0h�E`�B�HFR i���cC���f � 8��ԯ֯   ���.XBd���s
Pick? Press�v+=R�W�f�� ;/M//���/x�/ �/�/�/�/�/�/(?�Drop�/0/�? �?�?x?�?�?�?p/:? $O?0OZODOfO�OzO �O�O��Oi?�?,_>_ P__%_�_�_O�O�_ �O�_�_�_�_+oo'o�9oKo�O�uGRP ;2��{�jU^o8�o�o�p	 <�o�o To&T:L�t ������� � >�(�6�X���l����� �����܏	�0fX�����  ��  �S �� � �@E�2�\���>�HH��  �\�L��@u��iT^
>��P  D���Z_D�]�s>�N_�D�@
|�Z��ΕV��J� F�^_�ϔ5��*�k� N�`�����ů�������`��������t�P���菎��� �����ؿ��$�E���>�l�V�xϢ�s>��so^8	�  [��� ��F��d� ���-��oL�CFG ��k � ��g��P����o����	q	p,bk�K���q�x����� J�OG ;2��k
 l��s!��%�7�|�[��m� ������n������ !�3���E�i�{����� F����������� ASew��� ����+=O �a����b���//�mNET ��Vݑϳϵ�0&U�M_CHK  ��dc`��&E�LB�/ 
�&FO�BJ�/�(���/�'P�AIR�/ �&W�T?�$OTF 9��e�% D/Ԑs�=���A���b2�2��k ��P��[N�s_�? �?�?�?O!O�=�?�? OyO�O�O`O�O�O6O HO�O_-_?___u_ �_�O�O^_�_�_�_�_ �_)o;o�_�_o�o�o��ojo�o�ov/K�SE�TUP �V������5�KY`
 �	
��N/p/r/�� ^�r���������@��2�E�P`�o�����2m�����\`������\`F��
_τ�
�Z\`� ��\`פ��ˀ$\`����J�`	�
ׄ���u]P`�b �/�U+�+�/��� aP`��`2��P`6�`��.�z�es��Њ�=�`���ٛ��`� Q��`򀱖�`:�����n�ˀ"\`s��`��?\`�`������p�`���N�e������ m�`�����`#�F���+)����`%ˀ� �e0 &|�� Ȳ�`'���*�`(R\`��`�� Z�|��V��eP`��`+��fҀ��`��@���V�ïկ��� lj���3�U�W�� 7�a�C�e�������Ϳ �������!�K��� �Vό�2Ϙ����϶� ��
����@�"�4�F� X�rߔߖ�tϮ��ߚ� �����@�r�\�~� ������������&� ���8�:�X�z����� ��������1& XBd�D�~�� ��� $> `bl�����L/�o ���b �"WTPR 3��;
 �(/q�b�Me�v$2��/CmZa�ad �s"���(UaUa�(a�2�#h/z/�/9?�/�/ �/�/�/
??.?�?R? d?v?�?�?�?�?kO�? �?OO*O<ONO`O_ �O�O�O�O�O�O�O_ �_&_8_J_\_n_�_�_ ?o�_�_�_�_�_o"o 4o�oXojo|o�o�o�o �o�o��o0B Tf������{�G B_CHKCMB 2�S)ԁ!�q~�ROBOT �,�}X� Ҁy0��u \�2��q����r
���3�ƋҀzُ��� ��t���ɋ.�a�� |�����1�ğ֟�����|�DEBUG ���
����˯�����گ�'���L ����t�//��ELB���qn�"�̿ F�X�]�r����@�ӿ ���	��-ϙ�Q�c� uχ�߫Ͻ�N����� ��)�;���_�q߃� �ߧ߹�J������� %�7���[�m���� ��F��������!�3� ��W�i�{�������B���������FO�BJ 2����RрP��qM��7E`M�B��� ����@Rd9  8Y�{�}�� ������	/3/�*�
Pick Press'�������-g1�/ �/�/yC/-?/9?c?�M?o?�?�?�?�?Q+Dropc/�/�/8OJO \OO�O�O�O?�?�O �?�O_�O_7_!_C_ m_O,�_OrO�_�_�_ �_�_-o?o�O|_foX_ ro�o�o�o�o�o�o�o��o�_��GRP 2�����')M�	 <q�� �o����1��)� K�y�_���������� Ϗݏ��-��5�c�I�[�������0h�!n ��  ª�  �� ��  G�@�ٗ���}H��  �\�c�@�}(d^���  �J�ob�qs��PeD�@i��u���f�� of v�ܯ��ѯ��� �H�+�l�O�a��������Nh�������t����)Ϗ�5�_�E� gϕ�ϡ��������������I�e>�s�o8	�  ��}� ���Fzd�k f 4  TL_PRSNT_������ԙDHAND 2�\{
��Бfc��+�Mh�Z�=�O� ��s�������6�����=� �2�D�V� ��z�����������
� ���K.@Rd� ������ �Y<[`r�� ����&�
/ �J/�/n/�/�/�/�/ �/�/?"/4/??�/ X?�?|?�?�?�?�?�? �?)O0?B?OBOOfO �O�O�O�O�O�O�O�O 7_>OPO"___t_�_ �_�_�_�_o�_oEo L_^_0o�o$o�o�o�o �o�o�o Hoe lo>�~���� ��+�� �Vh��LCFG ���S  N��������ܫ���Ӱ<Ã�,���Ձ��xVr�ef�dӰr��[���OG 2�&�� l�ҳ!��S� e�w� �����J���͟ ߟ�����9�K�]� o��������ɯۯ�� ��#�5�G��Y�}� ������Z�ſ���� �ƿ1�U�g�yϋ�2� ���������Ϟ�	�-��?�Q���NET ���� 8�?�]ۏ�]���PAI�R 2��� ��H�P�P� P���U��*�<��� `�r�C���E�W����� ����"������j� |���Q�c�����9�K� ��0Bx� ����a�����,�߇�SETUP� ���P����K� 
 �	
zpƁ�߬߮߆�� ����/� /N/ o/F/h/j/������ˀ¾/�/�*2>�.  �� q_  �� F2�_42�Z� G���� ��0$T� 6�24��	>8)
&46���]ˀp�V���~4z8z8U���~4Q�aˀ��m��ˀ6�(�}1�1�8��0�=����4���90��A0 FJ��:D�4��0U"� s��?� ��:H� 0�p�RHA@A@��0��lF���m��1@E@��#X24�AM0)π��Y%0�0/�&�0UK����'�0���U*�(� ����b�A|�D�@����+0!0��΀@π��_$_6_DW l0ↂ/�/ �/d_�_�_�_�_�_�_ �_o=oo2odoNopo �o��[_�o�o�o�o 2'YCe�q �������o� C��?�Q�c�m����� ��͏�����?�)� K�u�+�e�������ɟ �՟��)��%�_��� S�u�������ݯ��ͯ �%��1�[�=�O�a� s���������ݿ���0�E�f�� P
� o�WTPR 3�z�
 �w�lm0�����Ϩ
dRR��LXؤ��D2ӷ����ψ��� �#�5�G�Y�k�}�*� �߳����������� 1�C�U�g�y���� \�������	��-�?� Q���u����������� ���);M_ q�0����� %�I[m ���b/���/�!+��C_3D_C�FG �NU����;"�"A�Z_CALIB [3��+��>�p`�b�P?a=,�/ �?n?�?�?�?�?�?O��?)O;O"O_O8&ROBOTjO|O-� ?.?@?�O@ORO#_
_ G_._k_}_d_�_�_�_ �_�_�_�G�_o;o�O �Obo�o�o�_�o�o�o �o�o�o70m T� o���Poro  �!�3��W�>�{�b� t�����Տ��Ώ�� /��S�N�w���� ���$���ܟ� �� O�6�s�Z�������ͯ \�گ�z�������]� �����z�����ۿ� Կ���5�G�.�k��� xϡ��*�������N� �1��U�<�yߋ�r� �ߖ��ߺ���	��� ?����f����߽� �����������M� 4�q�X�j���6���� T�v�%7��[B T�x����� �3E��R{�� ���(��� ///S/:/w/�/p/�/ �/�/�/r�/?�� @?a?s?�/�?~?�?�? �?�?�?O'OOKO2O oO�/jO�O�O.?P?�O �O_dO5__Y_k_R_ �_v_�_�_�_�_�_o �O1o,oUo�O�O|o�o �oo�o�o�o�o�o- Q8J�n�:o ���jo�o�o;�� �q�X���|���ˏ�� �֏�%��I��V� h����,�ٟ,��� ���3��W�i�P��� t���ï���v���� ����D�e�w�ʯ���� ��ѿ������+�� O�6�Hυ���ϻ�Z���$IC_AZ_�CONF ���������]�W��� ]���<]���MEM�BR 3��� �HROBOT��=����϶�}�_� �ߛ��ߧ�������� -�+�U�7�u�s��� ���������-�� M�K�u�W��������� ������%#M/ mk�w���� ��%ECmO����PROG 3��� �W�� �//$/Q/H/Z/�/ ~/�/�/�/�/�/�/? ? ?M?D?V?�?z?�?�?�?�?�?�SCH�ED 3���  �H]�����d]�
���Voxel Sched1Z�0OBOTOfE2oO�O�OB]N3�O�O"_]N4�O_j_]N5G_Y_�_]N!6�_�_�_]N7�_�_�Bo]N8o1o�o]N9Pgoyo�o�cI0�o �o�nnF $fF �FHZlfF�F�� �fFFV���fF�V  �2�D�fF�Vh�z��� fFf��ԏfFff�� 
��fF�f@�R�d��F �o��Ꟶ�?ٟ2��� �!�z�E��i�¯�� ���
�կ_���R�� ��A���e��⿭� 7�ѿ*�����r�m�3ǟaϺυ�������϶CFPACE ;3�� ����� 	 �D��  E	� D˻�[�B,@��C��[� �,�  ?�?aG�N��? |��f�xߊߜ߮��� }�������,�>�P� b�t��C�&������� ����_�:�L�	p� �������������| $6HZl�� �_����  2��hz��� �/���//./@/ R/d/v/3?�/�/�/�/ �/�/??Z?<?N?�? r?�?�?�?�?�?�O�? OO&O8OJO\OnO�O �OO_2_�O�O�O�O_ "_k_F_X_o|_�_�_ �_�_�_�_�o�oo0o BoTofoxo�o�o�ok �o�o�o,>�~-�LST 3�=�4�x{��?�l�c� u������������ 8��)�n�M�_�q��� ������˟ݟ��� @�7�I�[������֯ ��ǯ����B�!���DP_CONF ��=�����
��d� �px~5�E�pEz��p;� ?8Q�o@���]��`�q���o�SCHED �3�=�
��Deadlock� Prevent5� 8;�5�C�6� P�y�lφϯϢϼ��� ������(�>�D�u� p�z߫ߦ߰������ ���;�.�H�q�d�~� ������������  �6�<�m�h������ �t�������  6<mhr��� ����
3&@ i\v����� �/�/./4/e/`/ j/�/�/�/�/�/�/�/ ?+?����5??�?x? �?�?�?�?�?�?�?'O O4O]OPOjO�O�O�O �O�O�O�O�O#__(_ F_T_}_p_�_�_�_�_ �_�_�_oo,oUoHo bo�o~o�o�o�oF?X? �o(>Dup z������� �;�.�H�q�d�~��� ����ݏЏ��� � 6�<�m�h�r������� Ɵԟ���
�3�&�@� i��o�o`�Z�ï��Я ����/�"�<�e�X� r���������Ŀ��� ��+�&�0�N�\υ�x� �ϻϮ���������'� �4�]�P�jߓ߆ߠ� �߼��������� F�L�}�x����� ����� ��C�6�P� y�l������������� ��(>Dup z������ ;.Hqd~� �,�>�/�/7/ */D/m/`/z/�/�/�/ �/�/�/�/?3?.?8? V?d?�?�?�?�?�?�? �?�?O/O"O<OeOXO rO�O�O�O�O�O�O�O �O+_&_O_���_�_ �_�_�_�_�_�_oo "oKo>oXo�oto�o�o �o�o�o�o�o#0 FL}x���� ��� ��C�6�P� y�l����������X_ j_|_֏?�2�L�u�h� ��������Οԟ� � 
�;�6�@�^�l����� ��˯��د����7� *�D�m�`�z������� ƿ̿�����3�.�8� V�dύ� ����~��� ������*�S�F�`� ��|ߖ߿߲������� �+��8�N�T��� ������������ "�K�>�X���t����������������#����$IC_DP_S�ID 3�����V� � !gy ������	 5?lcu�� ����///1/ ;/h/_/q/�/�/�/�/ �/�/
???-?7?d? [?m?�?�?�?�?�?�? O�?O)O3O`OWOiO �O�O�O�O�O�O_�O _%_/_\_S_e_�_�_ �_�_�_�_�_�_o!o +oXoOoao�o�o�o�o �o�o�o�o'T K]������ ����#�P�G�Y� ��}�������ŏ�� ����L�C�U���y� ������������� �H�?�Q�~�u����� ���������D� ;�M�z�q��������� �ݿ�	��@�7�I� v�m�Ϭϣϵ����� ����<�3�E�r�i� {ߨߟ߱�������� �8�/�A�n�e�w�� ������������4� +�=�j�a�s������� ��������0'9 f]o����� ���,#5bY k������� �(//1/^/U/g/�/ �/�/�/�/�/�/�/$? ?-?Z?Q?c?�?�?�? �?�?�?�?�? OO)O VOMO_O�O�O�O�O�O �O�O�O__%_R_I_ [_�__�_�_�_�_�_��_oog�$IC�_DP_ZID �3����Ua�� d  +o!o�o�o�o�o�o�o �o�o�o"OFX �|������ ���K�B�T���x� ������������� �G�>�P�}�t����� ����������C� :�L�y�p��������� �ܯ���?�6�H� u�l�~��������ؿ ���;�2�D�q�h� zϧϞϰ������� � 
�7�.�@�m�d�vߣ� �߬����������3� *�<�i�`�r���� ���������/�&�8� e�\�n����������� ������+"4aX j���������'=jDL_C?PU_PCT84�B�  n @w��!VMIN_�]a =��G`G�NR_IOERR�  4[eDcIC�DBG �Ui�1-iicme�dbgD��$d�.�i�</,=�/iisv��/ /`/r!*/�/N/�/�ov/?�/�/
1�/k?��/D9)ud1:�u?�?=j�DEF c�Ue!�-�1��[0buf.tx�t�?y?�?�_BN�D_BOX 3�vUe� 8Ue�\OnO�42HCF��8�"1 %O4A�O�O�O_.
�O8_.dX`$;5"�D�ZSTATE 3]�GK �"'_ �^�_�_�_�_�_o.�_?o.ocoRo�ovo�o.�o�o�o�o�o#G.6wf������/K����&_-�_Q��pPS�I��
�(RNP�Tx�M_DO��"��uPL_SC[RN� �����TPMODNTO�L·��_PRTqY��n��VIS��ENB·�F��_�FFRCVR�x�I��G�M  R���b�D�RSMPR�GO���o�����$IOLNK 1���ߐ�0�B�T�f�x�|���MASTE��2��OSLAV�E �����_A�UTO�B��ܨUO�P����YCLE��ۤ�0_ASG +1�GI�G���n� ��������ȿڿ�����"�4�F�X���A�N�UM���
ݢI�PCH(��RTR�Y_CNb���O�ɂ_UPD���b� ݢ��B����@ߝ@VP_ME�MBERS 2�:GG  $tGU���"LtKW���V�RCA_ACC �3��K  T��� }�� �X +� 6+�h44�a��K� ���ߎ��]�4�ܕ�B�UF001 3���K= |�u;�L�(�} uB�pJ�} u5�t� �}@uC�F^.�}`u0�  u0}�V�*V��V��V�~Y�x�� v�@u1X�1~�U�~�u<6?�0~�uBV��`~�u<3�A�d~u�}� u���uG��U�� t( ���g�8  g8x��x�@��U�x]�xe�x��u6X�6x�u�5X�5y}�y��y���y`u7
Wjk�y]�ye�y����yu�z u�0u:�z u=[���z@u6g�8UzU�z]�ze�zm�z���{}�{��{���{`�{�uA�5A@ {�u1� e{��/L�E�{u�A�3`}|��Xi�|���|��|`uGr_��|�u5c��D|�uCuCG  |m�V��2 �^2�u;  <�u.�xD��L�`�XT��!`S�\�m���d�\�Hl�Bw�2pt�< 9{��CP1���B�21X��V��u<� �� I��u�V����� �������V�������<����`�@����/.F��V�p$�u0�h@�<�$�P@D� =fS�U�8\�V��d�9�;@l�u=<ku�f�@|���t(����ެ�H_���XP��fA��$��PX��b��x��V���]�q�� _������3)2�B�<�J" E�J"M�J"U�C ]�C  e�C m�C u� }�  �� �� g$��"�� �"���"�$������$ ���Ԃ����"�� �g$� w$�� �  -40�$4�40=�22 o$L�40U�40�$d�k m�r2u�r2g$�kw$ ��k���2�$�� ����2��2�$�� B����2�$�� ���2� �2 �2$�ԖA3��K 4��OI?�B��!�ѱ!�!�����HIS�� �ܳ� 2022�-04-1)2B�C �� ��� �D �D�"� i"� �"� �@+a: H  � 7 	
� �$ )X�a9 �`   ' $����@p�Dx �  % &�  �@c�N_`_<�T��`�HY"�HQ�(��;N@b�@ �+ �O�N�@��@�P
� 6S 
P�QPJ@�T%PQ-P� 5 5P Q���D� �@/ ��   . ��&T�&T�&T�&T��PjAT�ZKA�I+*�PH��2G�T�@�a�S�P�b��1  �RW��b�� , 	�@�!c�@�b
��b P�bP�b�аb%P�b�-P�b5P�b`07PP@!`�b)`�b1`�Qc9`U8P]A`/�@NI`�bQ` qOT�Z3 �L�b���b�_�V R�H(�o�o�i4ߐW-Pr(5P�R`.+`L!`�r()`rx-��KA`�b>I`3 	 UQ`�VT�Z2�L�b��U,�I�@%/P=�h|0RW�#  ;��*�A�@5f@X�@r�
�rPrP	���мqV�o�f r!`9��_)`�r1`�r9`�r�sT�Z�"�O�O��\�R��@��@rm�6�PZP�aQ����l�r��φ�rI`�rQ`&��?T�Zi"�� �_�JiB�@iB
�iBP iBRajA��jA%XiB5P iB`iB!`iB)`iB1o�CojA�I( �O�OG~dYtd��墍`���� W����墉td�@T�[�P7�@[PT�P�h�Yi�d%P(;PC�-P  35P" Pb�t���t_�_D᯶�^���q^�@�b�PxaGP0RP2T�0���P `%P��}`-P )  5P*đ@`$�<!`h��)`0r��d̈́d��d
��d�dYo���ؿP� ��td�tda�QdB���y�d��d`���dd��]�o�r5 �Ϣϴ�xb������ �x��#�d2ܰ�m�� m�ߵ�)���!¦ؤR ���֤RE��R��֤R �h	�?�u��I�[����c���ڨu����������`sɟ$�6�H� ��l��ߐ�����������I1 ��Ưۙ]�lA (�08@ ]U�lAH@P@X@U`@h@p@x@� ]�lD���\���� ]z���'�/�7T�?�C�K�SU�[�c�k�s��{�lA� ]�^lA� ]�lA�U����c�`	~�ۙX��X�YKAYn�#Y�+Y�3Ye�;Z	AFZiK�Z�SZV"` [mc[Lk[�s�[�{[�_#\#�g#\\o#\m�z \&"� aA�!-�$�"� �a�"[�ܘT�TM�T��3(�4w0 T^"8 Tf"o@ UCUMK�U�SU�"` U�h V�"p V�gsV�{VV"�� Wg#Wi�r Wmlw#W�#Wۇ#�X�#XR�#X�؟"7�ܘPDPw�P
2  Pf"({ P�"0 Q3�Q;QKCQ�zKQ�"X Q�[�RBh R�qnR�qsR�{R�"�l3�i!SFo#S~w#�S�#S�#T6�#T"�#TZ�"��ܘLIUSTT zTT(TT0 LJ3�Lo;L6BH Le�KM��VMG[�M]���M�kM�sN+{Nd_#Nޞ2� N�o#N��w#O7#OM�� O��"� O�#P	 �"��J_\_n]2b�P2bP�P2b�P2bP0dX0dU`0dh0dp0dx0dU�0d�0d�0d�0dU�0d�0d�0d�0d�`1c��I_CF�G 3�� H�
Cycle �Time�B�usy�Id9lr)tmi�!�=OqUpvq�Read$w�DowCx?_�Tq�sCountq	Num r*s�Q��}��q��SDT�_ISOLC  ��	�����r_�USEz@�{�J�23_DSP_E�NB!� 5�OBPROC>��OqM��G_GROUP �1��{�d8�?]�����E?��ݏ�Q� �*�<���`�r��������y�IN_�AUTOc�(�PO�SRE^�.�KAN?JI_MAS�@e��*�KARELMO�N ����y [�t����������2�v�b��P���ޥ��Q�KCL�_LԐN�1�$�KEYLOGGIN�P� ��,��p�LANGUAGE� �z���DEFAULT� ���LD�a�@�O�KyKx�u��G����E���>� .��� � J ��'�"g  ��t̬�MC:\RSCH\00J1D|e��N_DISP ��$�Ky���ƴOC+TO"0�D��r�AB��GBOOK' ����QOt�����PZ ������ ,�>�P�`ݚrOtr�N�	�Ŭ���QZ߿��F}��_BUFF� 1��{ ��jE������Iw 9�K�x�o����� ��������#�5�G��t�k�}���E�z�DC�S � =���oܹ����$�6H��IO 2��� � }� �p������� �!3EYi{ �������/�/1/\ER_ITM�~d���/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�?8�?��_"SEV�$�][&TYP�~y/�ZOlO~OM��RST�1���SCRN_F�L 2�j�p� ���O__(_:_L_^_F�OTPG��IB��NGNAM>�Kuz�nE�UPSM�GI�@��,��Q_LO{AD[�G %�Z%
PRT46[��1k_�MAINT�_�R?�Z  (% odoS�Ro�ovo �o�o�o�o�o�o- Q<u`��� ������;�&� _�J�����������ݏ ȏ��%�7�"�[�F� �j�����ǟ����� �!��E�0�i�T��������ï���*iXU�ALRM.��Q���"E���Q9`�T�P����P1aCP���j	~�����%mG�_G�RP 2�M� ���	�Q��P��P#�䵲�̿޿ �h��F�1�j�M�_� �ϋ��ϯ�������� 	�B�%�7�x�cߜ߇� ���ߵ��������� P�;�t�_������ ��������(��L�7� p���e�����������  ��$HZ=~ i�������  2VAz]o �����
/�./�/R/+gD_LDXDISA�P�[�A2`�EMO_AP�PE� ?�[
 �Z+�/�/�/�/�/?�?,?2`FRQ_C_FG Ǜ�X�[?�&�@�Ӣ@Ӡ<Z�d%/<�?D>���ț��R	 �16-AP�R-22 14:?24:30 Ӥ�<�31:12�?C8�:04OC9:3L)O�341'OUF2CI �?Ц�O�O�OB/ͩ�U��O�O�ET�s�.P�T�t�6P�T�u">PQ�L,�(HOME_I=O��C_R0��k_ӡVW_Tb_t_Z_�_ �_�_�_�_ooo(h �OpoWo�o{o�o�o���ISC 1ɝ+ �_��Y�'��O`K��oC_M?STR ʝ+�w�SCD 1˝-� x�t��:�%�^� I�[��������܏Ǐ  ���6�!�Z�E�~� i�����Ɵ��ß���  ��D�/�h�S�x��� ��¯���ѯ
���.� �+�d�O���s����� п�����*��N� 9�r�]ϖρϓ��Ϸ� �������8�#�H�n� Yߒ�}߶ߡ�������6�MKU1̲}�1��$MLTARM�T2��7;� ����0z��l MEgTPUy r3���y�NDSP_CMN�T��u0��p ΀�~��q�1����P/OSCF��3�#��RPM�� �STO�L 1ϝ+ 42#�
���ъ��� ���������������� 4(jL^����������S�ING_CHK � ��$MODAFS3�+�G;�B�DEV 	�*	�MC:�wIHS�IZEy-�@�FT�ASK %�*%�$1234567�89 ��DTR_IG 1��mlJU��?F/Y5/v/]�Y�P�U�tEEM_INF 1��;�`)AT&�FV0E0{/�-)��!E0V1&A�3&B1&D2&�S0&C1S0=>�-)ATZ�/F?-4HJ?r?1f/�?)8A�?�?�?�?�?O$O �/IO�/? ?2?�O V?�O�?�O�O�?!_�O E_W_>_{_.O@O�_dO vO�O�__�O/of_So o_�oDo�o�o�o�o �_�_�_�_�_ao ��o��no��� ��9��o�oo�"4 F��ɏ|�$��̏ �G��k�R�����T� şx��������ҏC� U���y�,���X���ӯ������ONITO�R��G ?�  � 	EXEC�1��:�2@�3@�4�@�5@�
 B�7@�8
@�9��;� ���?� ��K���W���c���o� ��{����������������2��2��2ĸ2�и2ܸ2�2��2� �2�2�3��3�3K�FR_GRP_SV 1��+� (��@+<5�?�Y>��o�9ȕ���Ǽ��{���_D���� �PL_NA_ME !_�7���!R-200�0iC/125L� Base G4� S��RR2�� �1�����07�Y�	X d �ߑߣߵ��������� �!�3�E�W�i�{�����������
�2 ��)�;�M�_�q�����������u<��� +=Oas�����p  ��\  � � ��  ��  A�  B� UT� �u
� �� ~@���  ��� �� B� z� � � CuCuP �E;� E@O D��=�D#�>>#JW�  6:gE�d��g�E(�}��Z����~��/��������/}��:.�h0�������#3�P�'{%���/�! �!�!�%�!{%�%�%�!@�!{%��)�%�!m8N��%�!�17�@�(J"G4�"7<�&� �)c?�{?�'72?�2���?�1�1�%�?��3�!�8��!�=چ�� !C#A�?!C��`IC3OFFp �EnB[OQC+DF �?�6��O�77�O�N�� EJH�E:�`�E�
� :� ��  � _.[�dS� K_]]A_�_�W�@
��]wS��W%��_�_�V  A��`��iep� �c�����&oc"oPoa�
?`�CdB@�oi��-���o�l`�f��/�y��`kbl6 ���� �@F5?� q���?� q�@�6�6�1�A~;�	}l#r	  p�� �,^���x�\p�� �� s � � ���r��K�l,K����K��2K�I+�KG0�K �U�\A�U,_��~��6@ t��@�X@I���r,p��S�N�����
���?������p/��}Ð��a��k��ôW��  �8��$ �������R���� D���W�ʍ�}������_!��U	'� � ?��I� �  ��Ca�Z:�È~c�È=���{��r@�������a��
��bvTʏ؏�yN[��  '#�<��$�?���r0���r8���B� b�C�X�Bg�
�� }��k�qt� �_cb�~-���u��BC`��[�ǥ�[ ��(q�R�_��_,� �P�;�M�@�`�P�������� ,� �� :/jdSD�?��ff�_��ӿe� �����q��0ϖ>�?Lb�qC�(� l�PuȐ��qkskt�Փ[�Dܮa;�x�5;��0;�i�;�du;�t�<!�ڣ���A�f�#r�c#r�?offf?��?&���d@��A=#3�@�o[;�˙ ���D�pus�w�� �Wt��߲������ ��3��W�i�T��˘��FР|���x���@d������A���E�PCҐ'A�Ь0��� |��������������� 3WB	ꟄH>���(��_�G���KG��]F����C��FmĤB�=( :L��?`�qO���c�����cA�РA�$C`Bb'/A��L/��Ū�?Ƀ�z/�/�/�/˙�mآ��n�/C���` Ca�/�
�$��� �!71�p�K����bC@_;CL�n�BA��Q�>V�^È�����Y�\���Q�?�p���Q��hQ��@�G�B=�
�?h�Ó?�`�����W���ɰ��B/
=�����Ɗ=;�K��=�J6XLI��H�Y
H}���A�1;�L��jLL�PBhH:��H�K�O@	b�L �2J���H��H+UZBu�/pO�?mO �O�O�O�O�O�O_�O "_H_3_l_W_�_{_�_ �_�_�_�_o�_2oo VoAozoeo�o�o�o�o �o�o�o@+= va������ ���<�'�`�K��� o�������ޏɏ�� &��J�5�Z���k���Ώ�Gϭ���� C�a$/؟ Ĉ�9����CVF��E�␘��;q�,0��yKr�u�� 
E��Н�c��� (��_3�hꯣ��������N����k!3�lC�7�I�W�����c�u��t�.3礁}����k����q'�3�JJ ���������C�1�Jl%P��PuΔ�������Ͽ�����A����>�)�N�{N�<]߄�  fUw�9� �߭�����
�σ=�+�a�O��g�q��̕��)Z����  ( 5� �����-��Q�?�u���  �2 E��k#Ew�L�����q�cB�! !�C�	08!  @���k$���0BTr#n���}��Ӥ^�0����?��k(Ec$�k �g$r+
 �0BT fx������`�//�:j"��_��u^3��$MR�_CABLE 2��_� �w4T��滺z/bɯ/ �	� SϏ#�/Y�_��/ ?????I?s?�?[? �??�?�?�?�?O;O �?OEOoO�OWO�O{O �O�O�O�O_7_�O\��f��/�_�_�_���z_�_�_ o��*�#o** S#OM ��`)�}��� &j}lv�%% 23456�78901`ore �]o�o�a����������
�g�-1980/0�ao 00:�b *����`Wg�TE�STFECSAL?GR  eg�
��id%t�a
1s����:"J|HZl~� 9UD1:\�maintena�nces.xml���   	�j  ��DEFAU�LT��S"GRP �2�Dj \ w����&�g�� �1st� mechani�cal chec-k���U�� _�f���`_
������xǏ؍.�H�`�=��controll#erM�_�q���Q_`�_a�s�M_�MD���"8����ǑΟ������E���+�|���J`C����ҟv������Я��D�V�Grea�se bal�qr busho�4�w�����r�������
��CF�geB�.�t�tery���p۱������	R�d�&�P8�JϬ��bôg���f���-���������������`�z�aúcabl��	�
�C�<��K�R���
���ώߠ߲���a@µ��κC����n����B�T�f����aO�verhau�� 7��� x�������"�4����� �/�a0���.����� W�iU������C����� y���asO�� Y�-?��' �G��i{ ���_���� ///}/�/k//u/�/ I/[/�/�/1?C??�HIST 2�%U��0�7pL�=���Ŀl�K�50� � -944.�5 hours _RUN 91��5 ���?�?�1���0���3�����n��L�MG-3823.2O��4A[�JO\O"N�1�!��OĬO&J�1ÿձ���FŬ�fN'�8i�H5526.0_ �0v�3��������P��}�H9060�O���0*߃�����25�R���{�f-114o05.4�_	X ���_�_%J�/Xo?o|o�z3SKCFMAPw  I5�0' ���q�o�e�ONREL.s4���ap�bEXCFENB�g
�c�e�a�FNC�o�dJOGOOVLI�@ud�3\Dp�bKEYwGu=Pu_PAN�hbr�^r�b�07|c{SF?SPDTYPx�e��cSIG(@�o�bTO1MOT9�a�b�_CE_GRP [1�I5�c\)2	�b7�I�0�m���\� ��T���x�������� -��Q��u���>��� b���៘�����;� �_�q�X���L���˯�����PD_T�HRSHD  �)1F@ zQZ_EDIܰr�gz3�TCOM_CFG 1�mul�~���� 
M�_ARC�_�b+F'xT_M�N_MODEv��yUAP_CP�L��
tNOCHE�CK ?�k wo *�<�N�`� rτϖϨϺ����������&�8�q;NO_?WAIT_L�wB���NUM_RSPACE�o�b���߷���$ODRDSP����vxOFFSET_CAR8������DIS����PEN_FILE�q���C���PTION_�IOXjqM�M_P�RG %��%$�*���)�WORK� ��	s �S0��*8)0�` �)2���b��ᠡ�&8��(8�4���R�G_DSBL  ��7�a��J�t8ORIENTTO�`f�C��p�aA ���UT_SIM_DRU��b�a"��V��?LCT �۱g�ad���`��_PEqXװ���RAT׷� du����UP� ����J0��AS9w�	�$P�ARAM2�����0��	X������ '9K]o� �������/#/5/&72�d/v/�/ �/�/�/�/�/�/?��<S/0?B?T?f?x?�? �?�?�?�?�?�?���`��`�,��  ���  ��  A��  B3@8�B��k#@H'@��  ��/@.@BJ3@z3@�v�u����P E;� EN"�D��xBMD^@�yEyB^@�N�A�  qEuB�DE��C�B�Ag�CE(��C�@�FZ��CJ@�F�H�B�AU/�G^"U2X�F�A��A�AR_�B�B.\u^�hkD�A�A��@���S3�P�W�U���_�Q �Q�Q�U�Q�U�U�U�Q@�Q�U�A�Y"e�Qms@N�@�U�Q�ENarA�A@�X�R�d�Rrl�V�D 2i�o�C�o�Wr@mBz@�b�� q�a�U�,s�Q�s@�A�Q*}چ�@� \s^q�o\s��`�snXvFp �E�@�r��sftF #v�A�wrA�$�@ ?ަ2@W�i������|���ȇ:�:��W%@���0�:���A���N���Z�J�p/@�W�����a�K�]���M��z��~�BJ@��"��������� O' 1��_,z팰`��l6��=��� @�e?.@R���?��R�t�D�a��ހ�;�	lb�	 � Z�� ��,^������� � s �� � ���"�H���9H�H���H`�H^yH�R���G�
��"�C��B�3@�@C4<�k�I����9G@z���k��y�º@n�R�d��v�#��$�{�Q����E�N� #�Z@ܿ��A��"���d	�����0��B��"�`��	'� �� ~�I� ��  �~��=���͢ϴ�N�@����˾���H��!N�	��Q�N��L߇  'X�d�/���B�*@>�y�:���q߃� >@  }�:�cb��-����O�B~��ւ���� ��"�E�G��k�V��z����5�������� �,�� :jA��>��?�ffُ �<��� ��F�X�b��8�o�}�?��I�^���(Ы�P��������Ӛ�A����;�x5;���0;�i;�d�u;�t�<!���.�Q��b���b��?fff?���?&\ �@���A#r@�o[zy���WM� R��P��@��1� �*N9r]� �����/�&/@���/�/(E�C��Dbq��o/�/ �/�/�/??<?'?9? r?]?�?�9)��=�?}� C/	Og/0O�?TOfOxO �O)z�&��GɑFO�O@BO_�O _9_�AQ�CA�TT~�}�f_C&_��_"X�?\?��ع_�_�_�_y��ض���noC�0���` Ca	o�:�T�x�P�Qva@I܊����bC@_;C�Ln�BA��Q�>V��������Y���\���
Yo����Q��hQ��@�G�B=ן
?h���oǐ���W�������B/
=�࿣��Ɗ=z�K��=�J6XL�I�H�Y
H}��A�1z��L�jL�LPBhH:���HK�J\p	b�L �2J���H��H+UZBuo��o ���	��-��Q� <�a���r�����Ϗ�� �ޏ���M�8�q� \���������ɟ�ڟ ���7�"�[�F��j� |�����ٯį���!� �1�W�B�{�f����� ÿ���ҿ���A� ,�e�Pω�tϙϿϪϜ����Gϭ���� �C�ac_� Ĉs��9�@�CVF��Ą����%{�߻`��K�ߴ�� 
E����ߢ�'���(���g_�h)�����Z��ųN��J�\�qQ�3lC�v����ⷢ��t�.�3��}����k����q'�3�JJ����:�(�^�L����p��UPP���1 �?��0�����7"��=D}h�{x����  fU� x�%I���?0|j��Ϧ�����)Z�/ ? ( 5�WP$/�/l/Z/�/~/�/�( ? 2 E�#AqS�E�L��&��q�qUB�`PSQ-�C�H``PqP@-�(?:?@L?^?p?�?�=�S@��?�?�?�?OqS?�C�X>UqP�Q9�T�[
 OoO �O�O�O�O�O�O�O�O�_#_5_G_Y_�j�R�����u^3��$�PARAM_ME�NU ?����  �DEFPULS���	WAITT�MOUT�[RC�V�_ SHE�LL_WRK.$�CUR_STYLv���\OPT1NoPTB'o!bC�_R_DECSN�P ��xlro�o�o�o�o�o �o&OJ\�n��QSSREL?_ID  �������uUSE_PR_OG %�Z%���sCCR�P�r����S�_HOST !�Z!�M��AT���i�0�B�k�|���_TIME�R��v ��PGDEB�UG�p�[�sGIN?P_FLMS��Ў���TR���PGA�*� ��?<�CH����TYPE�\�0������ 
�3�.�@�R�{�v��� ��ï��Я���� *�S�N�`�r������� ���޿��+�&�8��J�s���WORD �?	�[
 	�d��r�AL��U	JO>a��T�E����COL��o���o�TRACECTL 1����Q	 ��� �  � �]GA I@� ��!W�i�� �DT �Q�����9�D� � x����4�Ѥ�r�!��T���E@��ҽ��=@��9@��z����p a��Ub��c��d��e��Uf��g��h��i���j�ԋ�Ԍ��s� �]�]�]�]�����������a�9�]�0vo��� ��������������@������������	��Q
��L�������U��]�]�]� q�_��a��a��a��a��a���]�]�� _⦭Ԍ�Д� �М�Ф����д� ���ҩ��ҩ���$� ��,��4��<��D��L�иp����*��������ꀊ��H��I���P_⧪]�]�]�]䫨��a�d�k�s�*{�������a� ���a�$�a�,�a�4� a�<�a�D�a�L�4a�P<a�Da�]�]�]�0_�]�La�Ta�\a�]�]@�� ��������#5��PD��L��%��&��U'��(��)��-��U.��������U����������i �i $�i ,� i 4�i <�i D�i L� i "i <i Di D i Li Ti \i d i Li Ti \i ��i �i e$e$�e$ e$!e$"e#��$�$�$4�44L4T4R\4d2��/��0��e1��2�ѥ�q;� �0D��0L��0"�0< �0D�0D�0L�0T �0T�0L2�0T2�0\2 �0d2�0l2�0t2�04" �0<"�0D"�0L"�0T"��0*�4���0���05��46�47�48�4;��4<�4=�4>�4?�4@�4&`�2>`�2���2�����CP�BP�BP�BP9��EP ���EP���EP��� EP�#�EP�#EP�# EP�#"EP�#2EP �#BEP3REP3b EP$3rEP43�EPD3UK4S4[4c4uk4s4 #AT$AT4"EP<"EPD"EP@L"EPT"EP�BEP+AT!,AT\"EPd#�3EP �2EP�2EP�2EP��EP���EP S'T/T
7T?V:AT�BEP�B EP�BEP�BEP�BEP�B EP REPREPCAT�pCR��CRFATdEPlEPtEPJATREPSW MATNATOATDn�CRQAT+�CRSATT|EPUATVATWATUXATYATZAT[ATU\AT]AT^AT_AT`AT�EP�EP�EP �EP$�EP,�EP4�EP@<�EPD�EPL�EPkATUlATmATnAToATUpATqATrATsATUtATuATwATxATUyATzAT{AT|ATU}AT~ATAT�ATQ�Tr��odwdUd�d�d�dU�d�dc$�dU�d�d�d�d�F��0���0���0 ���0���0��0���0 ���0��0$��0,��04��l�s1��r1��|1��r1��r1��rk�a�$�a�,�a�4�@a�<�a�s�����u~d ɠT"ɠpra� �a�(� a�0�a��a��1�� 1���1���1���1��� 1��1���1���1�� 1�$�1�,�1�4�1�<� 1�D�1�L�1�"1�< 1�D1��#������ 1�L1�T1�\1�d 1�L1�T1�\1�� 1��1�L21�T21�\2 1�d21�l21�t21�Xb�1�`b1�hc� mĬ� ��� �� ô ˴ P���mĴ# �$ c� <"1�D"1�L"1�T"1� �B1��b1��b1�\"1� d"1��21��21��21� �21���1���1��B1� �B1��B1��B1�@R1� s����ƿع�Bɠ� ɠ|�ɠ�ɠ�ɠ�� ɠ�ɠ��ɠ��ɠ� ɠ$�ɠ,�ɠ4�ɠ<� ɠD�ɠL�ɠ"ɠ< ɠDɠLɠTɠ\ ɠ�ɠ�ɠL2ɠT2 ɠ\2ɠd2ɠl2ɠt2 ɠXbɠ`bɠ4"ɠ<" ɠD"ɯos1��B1��B 1��B1��B1��B1�Hr 1�R1�Xr1�`r1�hr 1���d1�l1�t1���r1�R1�Ss��{�������������$�$�k4s4Wd_d�gdodwdd.�d �e��U��r 1��r1��r1��sr߄� �ߨ��r�1�u�� �����) ;M_q���� ���//%/7/I/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�oM�q�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ����ϳo ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? ��C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/� A�S�e�w��������� я�����+�=�O� a�7?��������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q����������� ��%�7�I�[�m�� ����y��������� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_��_�_�_�W�$PG�TRACELEN�  ��  �_����	f�_UP �����8a@`$a�9`	a_CFG ��8e"c` 9`����qdo�g�ha�nMbDEFSP/D �Xl��`��	`H_CON?FIG �8e cW ����d�dM�b ���aPed�haq���	`IN~P`TRL �Xm�xa8�e+qPE�e��g�8aqd�a��iLIDQc�Xm	~�tGRP 1��i� ��B��  ���
��A�PH��@�r��ApD	�7 Ap�e	@�dha��y�zt� 	 ��ov,�(� ´# c�B�,�Bd��� j�T�����}�ڂ��}���BC5���.�� <�o S�3�l�/�i�����Ɵ ��K�՟�џ�D�/���pzi�r�`
 ��t @d�e@��F|mf��F_j(t�U�ʯ����ٯ���"�H�3�  �=�=�j O���K�������⿔f�)��)
V7.10beta1�f� @�{@�A&�H�qj�C`CְB�)��D1� ?�C���:Û� D�Q�A@ �qB ���p�q�C�q `� ?�I�w�C]�sŇ����pp�Ϳ�{�i��t�ۂ�����B���B�33C Y����k�B���������p���qB���{33B�ff�APlAN�WBZ���Կ�� пֆK�]�G߁�k�qc�A��*SYST�EM*��V8.3�382 ��5/9�/2018 A�e�P�׵��rS�V_T  P� $CUR_S�CRN`�GR�O3`&�PS_SAVE_DO`�;��E`$NO_R�ECOVERQ�R�ESULT:� �  
$PAY�LOAD`u�_UX}�Y}�Z}�I��uI��I��ARMy�1��2}�DO�aA�h�Q�MOV_PO�S��q�	����S�PEED_HIGuH`�LOW*�AC`%�=�5����.Q� ��M�q�� � $MA?X_PYLD�`���XISINERT?IA  �8�(��C��L�����?MOMENT���_n�SC���m�W4j�����IN��7 ��MN�����CL��PLD_M�ODE��DUMMWY11�`028��M,�s� � {$��_ENBQ��WK `S�ANG1L+��JAA}�JYBb|CC�D|��LST_t ��
$COMP_SW�`�}�XY4�~�Zp�� q� ��� ����}���ܳ���$I�`DI=S2� 8�X��S_G� | Q;���4�5�6����������1E� e�o �v��q�pyq�PMON_QUE��Lp$QCOU��,�QTHe�HOd��@ H��e�ISL#�UE+ 1��POtR`�q�$P) �BU� ,�\�RUN�_TO��dm DWATA�p�&�C��,��INDE�X�PROGRA������2��NE_sNO�$�%ITP�#�m INFO�	 �z �+�!��� ��! 2
 (��SL?EQ_NUM3 0�YP+?2�&�!SC�HKQa� 4�4 ENABw� P�TION[#e�ER�VE���9C# \3G�CFe1��$J� ~�"�$CA�R�8�?�7�`Z1_�EDIT� ��s�� K�93$H/IDE_��UGH�AUTW�ECOP�Y� 0LCc�MV¹0N:@>KD0�#PR�UT_ ABN�0O�UCHo��AP�_PRCREs��S�o6 �ME���IZG3� _RSET_DI�L� �?IN_FRO;3�A�D� �C�&DSP_qC oQTCH3`�p��-p��s�HS�TS� _SN���7�WRN_ALM_C�NU�DFi�_XRQ��JISq1' NTB��Q�E�R�P�C��P�RGADJ� �h�X_m�I�!�$� �V� �VW�XP��XR�X �P�NE�XT_CYC�Ce-L�QNSa5y�wQ�GO_]�$NY-Q�@EQW�@D6\a�F\�LA~CSa�Qp��@95�@ATEK#�]�IFY�&NAM�+ %�d_G~CS�TATU|~C'MAILTI�`+��a�EV�,�LAST��a*�.dEL�@f0� ��IhPEASI r19��FUr91D�Ev
�2O�A|0��~�Sb`��C!X���zrAB[!���E� 3�Vq�vB�ASP�vcp�sUPsD_� P�$�q�wRM>PRts~�k��s�SPK# q�t ��.d��	~Qr 2 �B ���6��r6��( @o���rb�ebAOP'DOU�#��I�Qu�PR^�f0/2GR�ID�![#BARS�86{@s3`�POT�O��� z!_"�d!�P݂��O� b4� � �� P�OR�#�l%�SReV�`)&��DIY��T_7 @�R�C \�3�Z�4Z�5Z�6Z�7�Z�8>���PF��q�!x $V�ALU�s.�7tp�|��b4| n5�R��!���a+�0AN-���aR�0E1+�?TOTAL_�dxp�B�PWIcI��W�R�EGENU�j��X��x�#E5z�& TR�s�BU�_S&R��j���3V�Q�4ڢ�2�rE��c��E!*�"&@�V_HƀDA&٠�GS_Y_���FS2 {AR&2 �BgIG_�@*�UP���e_� *����E�NHANC,! T �I�aG3��1P=�a F�#�p_OVRK#P ��B$�a&C����j2���86��ц�PSLG�Af0��7��E8��(?��`S���dDE=�U7�&|!�-Qe1�� !�B|EJx�W�eSIL_M|db��V�r�0� TQ�SH� �!�pC���V�ˍC��P_��P���M��V1 �V1�2��2�3�3�4�4��Y���C ؚ����IN��VIAB6 �������2��U2��3��3��4��4�ؽ�f��!�H�u��T $MC�_FI ^��L6�5ᑵ5�M���A���R�~� �\����KE�@HNADEDK�!��p��C���`��݁L�?���O !��D@J�,�㖷��REM�����a�C�����U�de��HPWD  ���SBMSK��COLLAB(�4�3���b0I=P�oN=OFCALn2�n� ,��FLt >�q$SYND���M� Co����UP�_DLYQx"DGELA���a�bY���AD&  \��QSKIPM i��� O� NT��h� P_� �"&�  ��P=�1K	^AK	s� J
��J
��J
��J
���J
��J
9�q�J2�R`� j3X�pT Vc��!���P�����!��t�RDC|���! � c@"�2R* +���R�A68C"59�RGE�0cs=��FLG !X�x�sSW�99�SPC�#�aUM_� ��2T�H2DR��  ?1  8���[0;11!" l~��0Pº�o3q�AT���C ���@D6"P0�$�[0�9���#��HOME�'" ��2�#���//%/7/ ��3�$Z/l/~/P�/�/�/�'4�%�/@�/�/??1?�'5��&T?f?x?�?�?�? +l�6�'�?�?p�?OO+O ��7�(NO`OrO�O�O��O L�8�)��O�O�O__%_ �D�SQ�O1* � lq��� i���E4d+�a��R8��SIO����YI�P�P��P�OWE��, 8�P��
 ,�2�� -��8b$DSAB5��`r1���C��� ��RS23�2�U. �.MU<��\�ICEU�r���E��PARIT��0�OPBy��F7LOWM�TR�P=�X��CU�`M4s�UXTAR����EORFAC�d��U,�� K SCH�z�/ t~�G��pE�C�$����OM$6�F�Af�IK��p�`�A��$`T�P-����. lxOs��EFAx�����RSMF��2�CK 0 L(J���7�7pM�wep�QEa�NE_T����D@�Y��s��(�uCTRL/_ 1 Gp�P2��A���FFi����q�PX�r�p�a@��GPM�c$SE�GFRA���=�c�M�G�q����u/20 *�P���r
� O,�TS��r�r��p�v���p�qDIOz�2 �����vU��vVz�3D �*�DS��+�kp��$�`_DR��n���A%�1�Vb��&�Y��O0��D%�2$ƞpAL��C�w�IN=F��_HAP��a4���YS�AJ�qe�����%��p�q˖5�I�TR�plRZ_OF�FT���PAUS_�������g�$MNT�qCM�p���Kp�q�q�4� Ӗq�ԕj��t��Іp���{�B�CHK���QUb�a����Va2COUQ�RE9G�t�ALA��`8䡍��SPG^�Va�A�f�FG���_�ebV��q#��TՓkq�aMO�#OU��STE��?��`S���DI�_m�ꦜ��[`OPT��UH��?���� ������֒7�ܚq?�{EC�Q5 8� ���#�sȠD��d�O`����V`�DI���{�6 D $UΊ�MSG�q��EV����ED��Dp�P��SHA�7 <���td��v�� �{`Ppq8�) W�OU+�A|�XZ6EEX pIO��qp �`���]b��d�ѶaF+�WRS�n_�ZDExO�E�VFRIE���qUg�M儌�TO;OL��MYHG��r�LENGTH_VTؤFIR ���P�c�q`��Ub�V_t� 5 �QRGI�ßWAITIF��X�#���G2�G1 ���/�@�Pt����O_,�{�t����`^������TC��8��Y����GM�rq9 @>�E�a8����/�
u��
ugt��}�+p��:X +�M�pC��q��1�E�e���G�W�/�E�+�Z�D��LO�J���  ��j�~��gX��� 29�JPI��O�1[��`2*M�2��3M�3[ڮ� \���!�V���Ц��$V����V�VDw �� ��u�p;,v��P�Ä��b�$z����lE½���=��T$���P!R���HSa fa��q�P����Q< 0N` ���:��j���;s��`�RQ  �
?@��S*a= E�xR-�M�o�>��4�N)`AX�a!�A�!�L�����THI̥p��LIuw�FEgREN2�IF簄CӌIM���V`G!1��O��A�; M&_J��%P��T	�RT�S>� ��`J�[p]�,�BD4�Cˣa z�U�����^�(��C �IN��W��Q$TBC[_P��CM�D�!jvLDR+p�Dq�!��������SWIT~jR%/t�R>�ATAq?܂� |�} >!$VALU1��P�&���@0b�! � 2? �SC�*bA	� �$ITP_��ĲJ�\3�TOT�\3�s6J�OGLI�cb�_PĂ��cO���.�AXtŰ�fK��MIR�1d�4Y�M��5AP&����E��jvűSYS��1��PGFBRK�u�kvNC�I�Q  ,B�7B^2V!!�\3�0BSO��\3�PINcE��6'a�V}����dcFSPD_O�VR��T��LD�B�3OR�GfP/��F�F��F�0OV�5S!F�J}�CM�F�FC��2]�X���bLCHDLY�7���D ��0aW ���WR�0RO�cxoA�0C�  @� ����ERd����0��WD.�PT�AoA�� �5�@���Y�Fp��4a!� ��Bʒ�]$Za� Va�Vq3�T30�Bٓ�FAMCa 0)p8ewRRo_M`�bx���s�PT$CA�0|���T$HBK[qPjv�aՁ��eIx�� PA�j�a�i�d�e�]e�a�SDVC_DB*�q?�G�pw�'t�1.zwc&u3.v}PADk�G����@UR�� �t��ABc�L�ڣ�u��1ha�0_AU�X$FSUBCPUG��pS��SK� d�`p���wH dFLA!yHW_C��V0������AC�T�$U�NIT@D:�3�A�TTRI'@G��pC3YC1��sCAsr�3�FLTR_2_F=I�TARTU  �2xtB"ҡTLP�;���CH_SCT�F��5�F_=�ƂO�F1S��b�8�CHQ���8���RSDF�� آe���`_T5hPRqO_p�S� EMP��04CT�O ��Xz�2�G%ERAOILACs��ME0LOS@��{D��~u��~twcPRp� �F�Cq =	vSFUNCR�RIN��$����!3RA�r� �`.�8�0�d.�WAR#�`#BL�E�_�AX�T�[�T�DA>@/���_�X�LD�p�@]���t128����TI�����T$�RIA,� #�AF�pP�A����oP���p�bO9I>��VDF_��rSKPD�Lܱ|�A]P/HRDY(�Oذ�!�԰Dӡ�`�MULS�E��'C�wa{�J�JJ�B�G�KFAN�T�MLV4S�WR	N絉�Dd��a�)7�;2$��DOWJP�p�ª6�STOS22E_KP�vAU`� |eZ�O_SBRr�gŀ0r�3�s���M/PINFvI��Ĝ����REG�+�D�G�b�VZ����qP���P�PG1B �] y�$6�$Z��C2-1H0C� ��3EG�j3�@F(�ARn0�s��2���7Յ�
EAXEv7R�OBs:y s6�!0B_��UCSY=@b�3@��S��WRI]P;���STRr5{`2@�@E"��0D���I�-P�B�ЃQ��
��c`O�TO��0�AR�Ys31⯑ct 1�1FYI@�3$� KO���Q�D_�ӃQtC�x�XYZ�:��5��OFF�PP�)x�l�5�Bq0�����*q4P����FI@����O�B�D���4�_J�12�BW%$h?�	��6�BUS%`�B'�_�C���6D�U��B�7TURB�X裘�?��X���`G�FLE 2P�s5�ȶ����8�B�Q +1B0K�pM�tB��9�u��w�SOR!QW��14���3�Cޠ @	 Q��f'C~1��N{OVE��M�� !�ÜӜқ� ��!����%���� ����0� /r!����%�%��1E)R�18�	ƒE]P� $ғcA8���&�`R�=砡�v��AX`S 2���!v�S���� ���������X��@������ �1�@ ������������ ���)��)��%)���5)��E)b!V)DEBU�$��z�1�Rt�AB���a�A|9V�`
� 
!27s =I5�qU7!�U7��U7 ��U7X�U7��U7��U7��d�����LA�B��G�sGR�O��G��|`B_ `�J�ԿC��o��62ApH.E]�:FAND ��pX}q}�[]�wG  |a��|�Hb��H�|��NT��q�SERsVE�@�D $���2�ACQ!�@PO �R��P+��A��B���E  $.�BTRQ��
�C��2PFW�2EU�~��_ G l�"a1�ERR�bI�`V���lQTOQ�� Lf����VR�eG�E%f�r��C"�QH ,�AU7P�F�RA�Q 2gG d�R�c��TnP I��$� �e�B�� ,�COC|��PJ  ^[�COUNT�� ���Sx��K/� �M�@�@�ELAY��MbVA��\Mb�qꡘf�9	yc��CSF����fK���b��d��d�ws�bV�g��cFX�g�wYzZyNUj4zV4zWuHP�` �c�frF�st�}wЀ}w�`}wp}w��S�FI0�jIG�DO�P0�Mb�q|D�sr4ZLb2QeL ��f�ߐ�NJ�`��*�S�F�Q�1+� �L`Z_N_CFGQM�S$�ƅ�T4�L@1ȩ�#�R�QP�\K�RdN �F0M����=	������F!A�����X��ڋഉ�Q<q��D$NuE��P�\�SS��DS� T O ̀F0SP�
�DU�K�����DI�����D�I���a�SEĮqZ�W+�;�_g$CDRwP��V����HELLP��P 5�B_wBASfSRSR�Ɗ}�|�S��ڡא1T�Wא2��3��4��U5��6��7��8�W.ʑROOea%V�{�NL�j�AB�Cn֒ACK26IN`T_CH:�j�?���-���_PU����OU�CPNw��*�𹑩V.��TPFWD_KARqQi�_QSRE�Dv�PM�N%�QUEᩐ� s�C=�I�53��y��8����y�SEMQ1}�r�]���STY��3SO�ti�DI���� �3E��l��PM�@���NRQֶy���y�$KEYSWIT�CH�/�����HE�s�BEATM0�PER�LEpR/A@.ȥU��Fl���S��D_O_HOMˀO�6��EFc PR������Ц�CH�O`sE�QOV_M9���p�IOCMe�U��� F�HK�Q# Dv�㧆�UXRC��M0��u f�FOR�C�WARI���qt��``�AR @4t�j�U��PAR���K�!�L�3J�4-A �8�S`O�L�0�S�R�UNLO4àVT��EDҠ' ?�SLCL��Q�Tl ���AN'CEL�B��I��t��DRY������WET�����_Q����)�<�հ�ZON1��G�?�2O�2?�3O�3�?�4O�4?�5O�5��ս1@������PU1R�p����SE�pt����RQ�9��W@P�&�^�U�Y%ABe����RSs �P�՝�:��UؐDEFN�� ��n�����������������=��6��6���7��7��8��8
��9��9��h��O�EN���
n��
 ��5�
��Q�
��m �
d��
���
� ��
���
����?GI_BCK�0���,%��(5%%��E@(U%M&�r&��O�����'�&Tf&�#�(��'�(SV��)�%Bk�H_R�C8�%?CLR_XF��(<'6YC,���K9�%�h<�%��O0L�&�5�7 I�7�<n��7�<���7��<��G�<��-G�%MAJ?��MFGG�3VG��3GF��SI�CGF��AUUG�D�J߰�J߰�J�BYV6�E�GT_N0�P�GS�%NO(ᇣ'Y�%POW`$�IW<�%�T_RD��iW �%򖠙%�U�%���W �\�6���V�6�VF -�V6FM�VdIg�\ �ig�\��g�\��g�\v6�O_�RI�e�g԰PLVu�V� )u#z�6')t�6C)t F_)t6F{)tRf� )trf�)t�f�)t�f��)tv6)0CKP8,�@�;�EQ_�K�c�;�FAU�d|�;�@��+疈;���Q1DK�����DA��م;����G����v(7z 5�ӯ� ��U �9B�  GROU�n�LAST_BIqT�Ъ�[ ERFJ�E0�G�_T֤���IN��葁���	I0���O0�p(��)V%�ƠSN3MT�ȑ�E_WIDT�6�7�SIZy�kPP�D�r�������T�P���м��	�FI�G]�0���0L��@��[ ��O���O�3Y��4��g�TO^� � 	��AIR��F�f�񒵣���KEF��P��~�ӥgTOG^�rCC%�r��G��^�SPXE������t�����5�	�6	�7	�8	�9 	�U���f���t����� ��I���V���c���p� ��}����I���� ��t�������I���V����c���p���}� ���.R��V  ��m���  �|��Ќ@SCFG��W_ � $��Dp����HAN��f���_wCTR�$ISe���T?�IE��PD���SA�ʝ�VO_�TYPE ��	�f�B�����a�"����/���/�I\�SMB_HDD~�� X v�BL�OB    ��SN�AS��Y� 0 $ADD�RES �$�$VAR_NA���%$M��PLY�_�zӉ�A�� Z� � $TIM�E��${�_Iޠ�	$�����Ҩ�CI<Ғ��FRIF��7 OSION���Us�=$֢INFO����BUS_ADR���2�-�P1TMS_��SPPTSK@�[ D �W!���$WLDR$XTRA_SH1P�J�$c�_MSK��CLj�X���S|��l�\ x ��NGLESTET�$DUMMYc��$SGL��TA���v�&����<����STMT����PSEG���BW�D���W�/��SkVC0@G?�] p��$PCS0NP>���	�$FBR2U�SPCT��U� ;�D@�R?�^� �$ހ�A00�З�1���2��3��4��5���6��7��8��9���A�� Ѡ�C��D���Ѡ�F��1��1���1��1��1��1���1��1��1	1�	1	1+	18	1�E	1R	1_	2��2���2��2��2��2���2��2��2	2�	2	2+	28	2�E	2R	2_	3��3���3��3��3��3���3��3��3	3�	3	3+	38	3�E	3R	3_	4��4���4��4��4��4���4��4��4	4�	4	4+	48	4�E	4R	4_	5��5���5��5��5��5���5��5��5	5�	5	5+	58	5�E	5R	5_	6��6���6��6��6��6���6��6��6	6�	6	6+	68	6�E	6R	6_	7��7���7��7��7��7���7��7��7	7�	7	7+	78	7�E	7R	7_ XF;�PR����l�_k�<`�� 
�;�(��k�`p�$TOR�АDtВ�1�I`&��EݠTcQ_CUR3REW�VaAX�������0�SYSLO~��a � �Հ0�c��"����$�c�VALU�eOP�(�$na�hF�aID�_L,��eH��fIN��FIx��+s�Ի$�� ��eS�AVk�b h 9$VpD�LCK�cr|��lxD_CPU|y@�|y���c-?t��a�TE����R c? � PW�� ��qL0��RXp���q��tRUN_FLG���	��tW���*����*��uH��K��t ?��TBC���� dX -$i�LENX�u�f�u��EL_R�,�$&�`W_|a�c1i�t2��MOtq�Л��ERTIAud#q؉�Idi��DE��֡LoACEMsgCC˃UbV��MA~���6��6�TCV=�^��TRQ]�~�t�u����Ѣ���J��Y�MDǔ�J�g�����
�u�2ǐ6����l����JK�VK���'��'��$JJ0l;�*�JJ2�JJ:�A��_�2�`�Z��_�*�}�N1����P�:��udLր�� !�d���e ``pGR�OU�`��.�a�NF�LI���REQUsIRc` �EBU���e�Ȗ$T"�2d�"�f��d��Њ�f \ $EN��^��APPR�C��~�`
$OPEN_�CLOSEn�-�)�������
d���g ��MC9�������'_MG&qɰC��WppӸȐ��ԷBRKҹ�NOL>�Դ��MO�_LI}���õJ!��Pb��2��:� �~�����6O���|R�J�  �d�>B�h� ������2���PATH ��������������'�9gi`>�SCAS��l`�ȱINh�UC܀�/�(�Cw�UM1�Y����7�qE*�S�2��S�:���PAYLO�A�J2L`R_AN6���L�p�ٚ���٪�ӵR_F2L3SHY���LO��'����5���5�ACRL�_lq%��!׆�3�H��`�b$HӲF�F�LEXb��d�J>h�i :u��� P�w�䊏4�P�������F1������Ə؏ ���� � �E*�<� N�`�r����������� ��ӓ��&۟�H�����TU��X�a ϑ�c�������)� ;�M�_�c�l�Z�~�����������b�Фj � ܯ� ��� `AT	��ƐELPw�]���J�i"�;JE��CTR!���TN:a��HAN/D_VB�bb��`n��k $i F2Ӷ؎�� �bSW�����d���l� $$M����^`ﱈ(�� �,���%=¶&Ap��öq�)̽Aݼ�`�A��A�� ޻�p�UD��D�P��G�p�t9ST�|1��|1N�DY�]�Ӷ�$�% ��j��׎����э��K��� �PW�`�i�`r�{ńōŖ�a$b���m ~ c�BxyF���AASYM���`���li`����_K��-�@�*��D@O(J�\�n߀ߒ�J���J���jS`Y���_V�I2#�X���PV_�UNI���T���J ��RE�R���T ��T f	�Ɛ�J�+�=�me�S�[� N���TCPPI�p Gn  �@O���P
����TCDELAY��� ��bSPEE>@� o X`p�dBU N]�� �b]���@�c^����by�ȐM%��$PRSq�f YP�E]��b_Фp |"� �bSE��¤�$�3p�WARNI��0EN2 ��OTF��qvv�_T��sM�AM�_tCc&�a_�HIST_BU__ q ,i P���PRy�q�f�rS;PD6tr ���g~* EARTBEהGSET�6p�CP��ARGM��FLGȕ�I���S��}�TR2Qb�BQp���{ぇ�]�REa����`��tOUTj�s p"�O�T=�Eˀ)q�F�IDl��j`U� ˱�(��c�% �St��d:�D�H�`Q�tH"tH��vI=�$DO=��  |�H�6su) � �"I�AA�s�����p�C��{��\��y�av � V`!ME_�sR�*�CT[�P��䒽����N�/P����T�NP¡ $DU�MMY1�$P�S_�RF��  t��@���FLAҠ��Z���GLB_T � wuu�i�U���F�!ʃ�w�`���ST�`�"�SBR\`M�21_V��T$S/V_ER��O"P��&ӣCL����Ax��`rA�D����x �ȐGTPSE�J�!�@�AD�b$FOR�C�BACK_FyI�/�BGLV#�A���CP�Ћ�SI�Zb�V�h�'��@ANAGE_ME$��$RECURS���$A��W� ��P1��/�  �D�GL�PEWj�y� 4�`��$�b$�Z�W�a��\#A\��1�  �ѳU׵�z i N�CPw$GI }$ױ y�ѳ
�j�G{ L�`,�!R}T�J"QE4�N�Y�N�yF{�V�TANC�_  ��JpR�!� |v�$JOgINT�a�  8ѳIM*�j�}�`*�Ea�y�S��@FĦj�_~� �U_�[?��LO>�O����sK�GLJ�Tp_sXMZ���EMP������KЍ��$U1Sڑذ��2z�
�Bo�{:�c �o�y��CEv=Ð� $Ke���Mi���ڰ�Ԥ��VEC��֨�IU�o�?qCHE>�TO�OL����V��REN��IS3���66���CH*��}��O�N��/�298���I�ق��@$RAIL__BOXE�a�oROBO@�?�ࡇHOWoq\�=�+�ROLMH���k(��p�����B O_F�?! �Ѳ�:9q��t����:9q���SLO����' ��Ʉ���k��y'����pIPA�NW ��M��Po�����OR&�������D��O�� �o D t�OB1 �Ђ�q�)�Qpq�!P��SYSq�ADR�,s[�TCH�  Q��rֈ��_,����tt��D�VWVA>�b� � �ײ�wu�pV_RT A�$EDIT#VS�HWR���B I9S}��INDϐ�)Y��D2Qg`4s {�+KE�a#�\�r�JMP��Lvu�h�TRA1�6t��y�ՉIJ�S�C�, NE���"'TI�CK���AM[q �d�HN��� 1@{��Xy_GWwD�΂�STYڂ)�LO���w��� t3 
�r,�%$,�u=�pS�P!$�Q ��ԑ酑��P�@XvgSQUe���LOꂖ�QTE0�P�RаS6t� 3�����""D���upT��lp�O�ݓ��i�,���<�pCH�?"{rUTsPU�QO%_DO�����XS��KvvAXiIn ��t�UR������$Tf����@�FREQ_�Ю�EET�"PҊ�EmAF�Gn[���CP0��>�8㉐ ���z�RkD�l� z���2���1P2%:�1B7>Vp)6�2Y8A�0Щ�&7�y<Ak@AV@Cp522�:D1�8D�>Df��<D�=�B�9CO��=C�=_,_>_PTa�$�SCw� � h�DS<�/�c�X�FAT�0Z1.�Ɂ��,�ADDRESz��B. SHIF$�^f�_2CH����I���A�TV��I�����rJ��A胇 
�I�
�bV�_!
�� \��"��m\!��ZRC�3"�",Z!��٢ZQ�TXSCR�EEs�T��T�INA��:��T,�p�a�!�B�`� T� ֠(u�R���V|!��|"|(t* RROR_����b�R�� ��UE6t� �,0��N������RS�U`wuU�NEX�vvdaH�S_Äf#ta�i�g#�!C
�`b�T 2m��PUE3���x��fqMTN_Z��r�� O��@�B�BL_-�W�
��S �m$rO��0rcLE�B;se�TO���$qRIGHDsBRyD��ACKGR��luTEX� muhqWID\�.�O �t,�[����C�UI��N�Ha � 8 $�pT_r�B�r�ϐRT �8㾷7����rO�A
��$�epUPp�RҐ��LUM��&�@ERV#��qP��@	���Ɛ� GEUR�D�F� ��){ LP$k��"E�aA)��qA����A�����5��6
��7��8x��#: P�nT.���S�����qUSR״'� <��ΐU0�S�0�FOC��2�PR�I�!m7�!j�TR�IPI�m�UN+DO��'����}�w�|�\�fҭ �� ��r5�>!G �zT��OA�A��O	Sm�֖R�  b���т	��������1 %x��Us�	����p�cs����OFF?Ъ
��y�.�O�� G1��v����ࠧGUN�u��� B�_SUB1��`SRT��4������#OR-���RAU�#0��T���VC�Cf`�� ��C?36MFB1t$α�VCR0Lĝx C�r�	�l���C��C\�n�DRI5V1&�!_V*���� ��D�MY_UBY�v�t����P�`���	��P_Sh���LU+BM7q�$� DEY?E�Xp8c	!� _MUb� X7qS�y`US�б���,bZ�G|PPAgCIN��RGa  |œ�d���#��¬cU��RE�r�A������S��� О<�TAReG��PO��� �S�9R���� d�}!d�qբ	T�l!RE_ÛSW��_A����$T�= O+��AA�@Mӊ*2E U`1���[ �S�HKe��e��!1J��P��E9A� ��WOR�pM�{ @S�MRCV�aW� �d�OqM�p�C�S	��v�����REFw������<�U� �#$�:���5���5��8W��֌�_RC�ۍ���J�S�K�³���s�S��d� �B�[��u��G�ǵ��RO�U/�¶v� ���PA2��`�PpP�> � ��CPA�Kn� SUL��E�3COX`T �E�4� ^�Pw�l���q��"���@�L����	ê��q̶�"��f���Gt +�C�!r@ �CoCACH�LO)���F�	�q�@�C�_LIMI�CFR�AT�0C��$HO��p� COMM��`bONpy��@g���VP��6�_S�Z3���6���1�2���w��O �W�ARMPFAIjO G�� AD5�U�IMRE��U_�$&GPf`;�!0P�A�SYNBUFP�V�RTD��esOML�@D_^��W#��P&@ETU4�/ Q�j�wECCU��V�EM�����OVI3RC5�VT< t%�$"f��"�_DEcLA��nQ'&.�����d�?aU�CKLA%Sã	��w0Gb�@I���/SWN�$�VLEXE3����S%�M��AO�FeLipI<�yFI� �'i��(+ē�O�w�K!� �§A��*���p"���n�;pORD^�A�9Q\�Qp��P��P�<�Tz��b�O��p#��V�B����`�E�R`�F�URO�7�_RC�Q�4 H�y�5���!�3�O  z�;A<�BFCT'0CF'SCO�2FCC�p}� ��{Ơ�LG��ZF��gG ��uHf�x����r�r���EzpAM!P%R���0M�����$�$gADJp0K����U����7ʑLI�N{�``��P5�� =x��MSPD�p&�"aR���Y �`I�"a'LNTjc"aM(0�ax�U�u@_ACCr�R-V���pZAB�C⥭<��R@3�
  T�ZIP��}���DBGLV��L�T� x��ZMPCF⥯ � ��K`{d]bѱLNKr
|JaI�㤇� �d��'%X�M�CM��C�CAR�T_�a_�P�P'$J�c�dD��b��b�g���e��a�UX9W�beUXEZ�vq�e�d�e*qq"y|q2vI\�Z!eO� ([�W�^ruYgPD�� ���:�6|�IGH~Í8#?(<�gV�;�_p>�� � �4
�`$B@�KKǨ�K�_�2~�,WRV	 F8@��3OVCP��b@�aS��0���0�
���IF��DV�TRA�CE��VY��^qS�PHER�� �� ,<�x��y���$PLID_KN�O7� N�̓��́��SV � ����=׀�ͅ`�̈́��1�C�  A	�j�U�����d��h����݃Mo! 1��\숌 �B�}�̓?���w����s��� I'�$ͅ@�̀ 5�=�9��K� ������ 1�ȝTͅA�  cB���ڑ̀C̀�B�����������:P�`1 1�����`4XL� Tool On�ly̓B���?��O�   A����G�� H�"o H��Ђ ��& Part���  ?G���ff�G�A IY�iI�@.�� BA����T�.� HT�]�Ht#�0��5� B�|��T���� H��H���G�d�Mi�[����q��F�8 H� H*r���д���|��G)�� HW� Hq]~-�M Dbl��Bb�̀��$� H� H�����8�&>�s��ff�Nƨ$���݁@H[��ɳS9�X|��S�y��G H4 HI�-����vƄ�Ȕ �0�� H�E�H�)o��ߧ2������'��<'�F��3 �#�5�G�ߧ4d�v��ߚ�ߧ5�������߂ߧ6
��.�@�ߧ7 ]�o���ߧ8����x����ߧMAD x ����OVLD  �������ث6�lQ z�吙��ծSCHU� c�
���lQ��׃UPD`����R\ߢ_C_`f
 ���'Յ�n�pCHK|��Պ�y�xAˏ݂a��_����`��� Ap��8�'�N@�E�Fw�)Zbi�� 9�w|����� ��+//O/B/s/'�8Y`�/}/0c� �/�/�//���/�/�/ /	�?4?9?/\�T? s?x?/���?�?�?/���?�?�?/V 1��сԑ�^����THR_IN��@��"deFMA�SSrO Z�GMN�qO�CMON_QU?EUE �Ն�� �� �Ns U�N�F��@END8�AYEXE"_U BE!P_�C�s�G�!�@��RAM %�J%�@0O��7R�TASK:�d_݁O#` �O��o��_ODATA��k���n��2 �uspv �swuj`�vgbkharck?vsm�o�o֮ek�axo`k\da  "�d��$�`�m�cX�ov��e�a�a��8r�ߐ ������>rb�� ��`P�`cuu^r���QINFO��	Km�������	� �-�?�Q�c�u����� ����Ϗ����)��;�6gI�t
Kl �f)�Q K_ahi�~~�Ga2��� P(O�=����ϟ��M� ��M�M�TDy�_EDIT o�9�2O�pWERFL�CXXCܣRCREP� �� B��FTТ�k���o�ʯFS`�ѯ��RGA_DJ (�A���?FP"�yA���A���=�~�B'&��FT��<���?%DIA4|��K�f,i"6�[�2y���r	H�@l[��BKA�UU�@e��*�/� **:��ƷCj�"@�FPꪪ�P��������kώ�D��	��!P ��[��8���:\φ��Ϯ��46#��z�����8�"@A����ϼA�f�C;�� ���;��O@(�R߷߲��p֗����@�8���@���r����\�j�N� �FP!�99h�^�A"@\���8�2��|�`�r� ������������� �R�8�J�\�n����� ��������W*" 4F��|��� /���n Tfx�/��� ��s/F/,/>/P/b/ �/�/�/�/�/�/K?? ??(?:?�?�?p?�?�?�?#O�? 	 ��1LO&LIO[OmDB��!��AƠB'��e�8��BF����b�t�$ �EpAJ�\���O\�dM&O�Om���Q6�PREF �D�P`b�SR?IORITY�Wf}�z�MPDSP�Qh�bWUT�V�a�q�RODUCT�Qe(�_��OG[��_TGe��R,��RTOENT 1(�� (!AF_�INE�Po)g!�tc�BoQk!�ud@oyn!�icmhoL��QXY�=��[  ;� )�� ��o�oP� �o�eD+hO a����������@�R�*�S=��+] %HOME�_IO 2 C_�R02�o�� =��j<�
o?�f���2022/�04/16 14?:42:34n���_T��������p��d��n�,  �:PA�MXm���SLKS�F�A�ެ�m�B��}�D�T�uQg��ENHANCE �D���j�A%�%!Oן�i#T+_=T�U�PORT_NUMԍSK�YUz�_C�ART� ¶�YSoKSTA�W R��LGS`�l��U�SUnothingޟ��ɯۯ�[�{�TEMP ��i�����_a_?seiban�OJ� �OZ���k�����ȿ�� �׿����F�1�j� Uώ�yϲϝ������� ���0��T�?�x�c� u߮ߙ��߽������ �*�P�;�t�_��� �����������:�>�VERSIkP�W�k� dis�abledE�SA�VE �j	2600H72��	-���!Ɵ����zo��� 	#�ROULSei������
���	����_��P 1�k��L��7Vh�7^PURGE��B�P�oVYU�WF�DO�V��{VW`��1��WRUP_DEL�AY J��R_HOT %@F�Qş5/�R_NORMAL(�b$/y/H'SEMIX/~/�/�QQSKIP4��Ex+�?'�&?8? J?�M�?{?i?�?�?�? �?�?�?�?O/OAOO eOSO�O�O�OsO�O�O �O__+_�OO_=___ �_�_�_o_�_�_�_o o�_%oKo9ooo�o�o�%�$RBTIF��N�RCVTMO�Uc�Q���`D�CR4!�) ��17�K�E?J+�B�X?4��#G�R��u�*+����[?]  ;��x5;��0;��i;�du;�?t�<!��o*�8Y��} �� ��/�A�S�e�w���𛏭����%RDIO_TYPE  S�=�ɏEFPOS�1 1"J�
 x�Home P?ositio8����w�%��q@+<6�?�[>��r�9ȕ���？�6L}<���5���5?�  ���$Ref/_Pounc9�#���S��ae�r������3���ПY���(����4���H�ѯPl�~�����5������I�������s�Ù�@8���\�n�����7������9�Կ�����8���(ϱ�L�^�pϲ�9�����)�������-��10���ߡ��<�N����2 1#�2����S�g7�����_��3 1$ ��,��&���J���n�S4 1�+�����\���}����5 1&�V�>�P���t�>��S6 1'����������	�-S7 1(D�hz ��A�S8 1) ���3�W�SMASK 1*�� 0�/"&�XN�O�&K�c.�MO�TE�`#�u(_CF�G +�.���P?L_RANG!�o��!OWER ,�Ye� �&SM_DRYPRG ��%�(?�%TART� -�.6:UME_PRO??�?��_EXEC_EN�B  �u�iGS�PDk0�0�8�a�6T3DB�?�:RM�?�8�IA_OPTIO�N�fp�'INGoVERS5A#���?�I_AIoRPUR�  G/\�O
�MT_�T� ��/�aOBOT_I/SOLCD.�B�ռӅ�BNAMEYL��iO\_ORD_N_UM ?�(�A�H72��n����xSLxRw xR�K�xR� G�S}�S��`PC_TIM�E�g�ix�`S23�2�"1.�iQL�TEACH PENDAN�`�c(��}��Mai�ntena-�CoCns�qo�"$o�f�No Use �~Uooyo�o�o�o�oׁ�RNPOE0�RO��CE�QCH_Lfn0/�N�	Cq~!UD1:izR�VAILYQ�9E�)SMFS�T_CTRL 2}1\J D%� ����(��OK�:�>o� ��! ��������Ϗ��� ���:�	�^�Q��� q���u��՟���� �/�A��Q�~�M��� ��Ư��꯹�S��+� =�O�a�s���[���¿ ���ٯ
���.����� ]�oρϓϥϷ��ϟ� ٿ�տ*��N�=�r� A��ϡ߳��������� ����J��n�aߒ� ���������	�� -�?�Q�'�a��]�� ����������c�); M_q��k���� �����	>� m������ �/�:/-^/M/�/ Q��/�/�/�/�/? ?�-/Z?)/~?q/�? �?�?�//?�?OO+O =OOOaO7?q?�Om?�O �?�O�O
_�?sO9_K_ ]_o_�_�_�_{O�O�_ �Oo�O*ooNo_�_ }o�o�o�o�o�o�o�_ �_&�_J=on]� ao�o����	�� -�=j�9����� ��֏�?���)�;� M�_�q�G�����}�ҟ ŏ����鏃�I�[� m����������ş� ���	�:�)�^�-�ǯ ������ÿտ���ϯ 	�6��Z�M�~�mϢ� q����������+� =��M�z�IϞߑ��� ���ߵ�O��'�9�K� ]�o��Wߑ߾���� �����*��ߓ�Y�k� }������������� ��&�J9n=��� ������	�� Fj]�}� ���//)/;/ M/#]�/Y�/��/ �/�/�_/%?7?I?[? m??�?g/�/�?�/�? �/OO:O	?�?iO{O �O�O�O�O�O�?�?_ �?6_)OZ_I_~_MO�O �_�_�_�_�_oo�O )_Vo%_zom_�o�o�o �_+o�o'9K ]3omo�io��o� ���oo5�G�Y�k� }�����w�ޏ�� �&��J����y��� ������ӟ埻���"� �F�9�j�Y���]��� ��ϯ����)��� 9�f�5���}�����ҿ ��;���%�7�I�[� m�C�}���y������� �����E�W�i�{���ߟ߱߇��$RS�MFST_SV �3������������*
�$�#��&�T������G����o�6���MASH_ENB  ��� ��PRG_AL_RM  ��
�x��é�DSBL��@�����4��8�@�5�S�5�
H�4�y��~�S���l���_CHECK 5!�>��MNCON?������DIALM 26��5�M�,	,\>��RUN��M��� SHARED ;27�� ����������	~TR�Bg��PACE1w 28�� ��@m�S������?8�?���� ������/'< N`r /���/�/ �/�?�)����=</ N/`/r/�/�/�/�?�? �?�/O�?O8/J?\? n?O�?�?�O�O�O�O �O�O_4OFOXOjO|O *_�O�O�O�_�_�_�_ �_0_B_T_f_x_&o�_ �_�oo�o�o�o,o >oPoboto"�o�o� ���o���:L ^p�����ɏ�� ޏ����6�H�Z�l� ~����������ڟ�� ҟ�2�D�V�h�z�(� ��������֯��	���2(:L�^� p������ſ濩�����1�6�3E�W�i� {���;ϱ�ӿ����� �9� �N�6�4b�t� �ϘϪ�X������� �@��5�V�=�k�6�5� �ߣߵ���u������=� �R�s�Z���6�6 �����������*� 9Zo�w�6�7���������% GVw:����6�8���� Bds/�/W/�/�/�/��/6�G <�� �/4�
<0 +?  �\?n?�? �?�?�?�?33(�=/ �/O�/FO4�d\@A? S?�O�O�O�O�O�O�O �?�?N�J5_G[d_WO iO�O�_�_�_�_�_o �O__/_Q_co�ow_ �_o�o�o�o�o#�o+o=oOoqo� `�/ @4��u$O ��o�i�2u�� +�1��>������� f���ڏ쏶���ҏ� F���,�^�����П �������֟���$��f�(�6|
���6�_MODE  �^ѩS =���`^zG/��a����	�����CWOR�K_AD�O��Y�R  �� �����_INT�VAL�($��R_OPTION�� �v�TCFB0>����!N����K�V_DATA_?GRP 2@<x!D�`P���ϓ��� �ɔ���;�)�_�M� ��qߓߕߧ������ ��%��I�7�Y��m� �������������� �E�3�i�W���{��� ����������/ SAcew��� ���)O= sa������ �//9/'/]/K/�/�o/�/�/�/�/1�$�SAF_DO_PULS̰0�a^�1�� CAN_TIM�ࡲeD�1R �A���������
N4	@}�V�c3*�U1�c �� �?�?�?�?�?�?v?O�O/OAOSOeO,� *�cY�2�DdR4U1H�A�A�Er4�m�p g�+��O�O��U1 _+W�PU2"�_  B��T��+_h_z_�_~�YT D���_ �_�_�_�_
oo.o@o Rodovo�o�o�o�o�op�o_:��L�kC

_Bwc3���;�o��'�p��m
�u��D�k�e1Gz� � �Y�*�eqe1Aa1 M1�����*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���"�4�F�X�j�|���������Oɯۯ� ���#�5�G�Y���|E ��������Ϳ߿�� �'�,�i���0�B�s U�}xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H���l�~����� ����������y�2 DVhz����l-ϳq��@�� %� � � ��pA (:LZk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�?�?�7��hw�P�? O)O;OMO_OqO�O�O �O�O�O�O�O__%_�7_EZON_{_�V����rt_J}	�12345678��rh!B!+̺�X@p�_ �_o!o3oEoWoio{o �aO�o�o�o�o�o�o "4FXj|� ����}�o�
�� .�@�R�d�v����������Џ�����BH)�Q�c�u����� ����ϟ����)��;�M�_�q��{;�j}�����˯ݯ�� �%�7�I�[�m����0����ǿ�yD�ѿ�� ��/�A�S�e�wω� �ϭϿ��������� �=�O�a�s߅ߗߩ� ����������'�9� K�]�o�.ߓ����� �������#�5�G�Y� k�}������������� ��1CUgy �������	�4�P8J/���v���YC?�A}��:   ��8u2�2�P} ��
��  	��226///A/S/b+K7��?d��P�1�3 4 5 6b/�/�/�/�/?? +?=?O?a?s?�?�?�?@�?�?�?�?O�.P&B(,B2ODOVOhOzO�O �O�O�O�O�O�O
__ ._@_R_d_v_�_�_���$SCR_GR�P 1C�|���~�Pt ��� �	 ��Q� �R�R�Te��
i�W� g.ooUo����RbD�` D��@�-�S�gRk�,�R-2000iC�/125L-IF/ 890 �e �RC2L 67�8�
V10.'03 p#h�Ra}!��*s�Qef�Q 2c�Q�#�QRa�Z&a8y	������~���H��P�jt�WBu�����D��sD����C3�@A���C/O�QC�L7A�jPAx�k<�&�ٿ������ � ?������oD��D����P/�Qo��Moк�����hp�T��~�#eBǙ��B�  B�33�B�	�����QA��+�  �aC��Q@9�A�T� ?�i����{�1��QF@ F�`������ҟ�� ����,��P�;�t� i��as�����������B�ίc����8� #�\�G�Y���}����� ڿſ���/�|c>o,�Q���Nσ�V�l�@��:���ϝ�O��`��	����1o2345�`90��e�5��AX�)�<� l�$c�PIЏ!=��A _߆ߘߦ�t��� ���ߨ�%O�!�1�P�EL_DEFAU�LT  <t����TF�HOOTSTRO�v�C��MIPOWERF�L  �[��W7FDOP� [�B��RVENT 1D����pz� L�!DUM_EI�P1����j!AF_INEO���O!FT��C�
�bg�!�R����V����!RPC_M'AIN���������N��VIS��������K!TP> PU�B��d:�!
P�MON_PROX	Y� �e��^����f�/!RD�M_SRV0��g{!R�ė��Yhj�!
��M����i�/!RL�SYN�`//:'8|/_/!ROS���,�4N/�/!
C}E` MTCOM�/� �k�/�/!	�"C'ONS�/��l�/C?�!�"WASRCdJ �m2?�?!�"'USB�?��n~?�? z��?>�?�?(OMOO�qO8O�O\O�O=�RV�ICE_KL ?�%�� (%S?VCPRG1�OZ"�E2__�@30_5_"�@4X_]_�@5�_�_"�@6�_�_�@7�_�_��@�do\9 o%k �D�Mo�A�Ouo�A"_ �o�AJ_�o�Ar_�o�A �_�A�_=�A�_e �Ao��A:o�Qco �Q�o�Q�o-�Q �oU�Q}�Q+�� QS͏Q{��Q� �Q�E�GQ��O�B �@�O�@��՟Qٟ�� �!��E�0�i�T��� ����ï���ү��� /��A�e�P���t��� ��ѿ������+�� O�:�s�^ϗςϩ��� ������� �9�$�]� o�Zߓ�~߷ߢ����߀�����5� �Y��J_�DEV ����MC:a���s�GRP 2�H��p��@bx 	� 
 ,���  +  UUp�p�,p�p�Up�p���c��+ p�p����(�a�������p�	�����
�虑Z� �,����������������Z�����p�����������XaH��G  �  U��`p�@p�#p�Ȼ������  "p�/�~������ ��0�������	 I���w^�|������h%/|
	_L  ���.p����)������*/�����/V	 �/f#�/�/ �V�5? �Y?@?}?d?v?�?
/X�?./��S �p����?��*?O�5 �eO�/�OpO��O�O O�O�O_�O`OE_ _�i_P_�?�_~��U � p��p�Y3� R�.���:fxO�_  o�6_,o^_{obo�o �o�/�o�o�o�o/؆_S�_ ��r
p�p��w(��~!,���P �p����
��?o��q�i J�K>i�o]�D��O ������ۏ�D� �>4�F�яj�Q����� ��ğ���ϟ��� B�)�R�x�_������� ү)������,��P� 7�t���m�����ο� ǿ��(��!�^�E� ��ٯwϸ�o������� ���6��F�l�Sߐ� wߴ��߭������ ���D��d �T���6�5���H�=?��%�?���::T�:�=�+N�N�l�<��>�����AS�X?���پ�">������C�@��&��Fo���d�����,I"��@����A�����@O�/��V!��%J�OGGING TA70 0�����c��g����?��29R�p9�{������[��k�`�ࠁ_A�V��?������v>o"[�����@�8��F�:X�d������o[�?A����N�A������!�@@�P��"�[��%��/��g�� �?7�G͛�9UU�k�������AT���?l𾅖�>�D�v���@��H��F�d��ߣ����[�=���
�!A���b���n@7؟d�a�&����Cq1����,��X2g���k῀h���!�@�?���:I�o�C �������ۂA�",���@�&v?���s[��� ��M�H@��C���e�£��C�T_Z�@?�����>&?<͠���-K@}�@�p��
	PRT50DROP ����=T��+g�=��=�,�>��Nl�H�N>�T�*�[����A�%�A�.墿���@��[�B��a��i*�Aq��B��n«V��Ac[��9���ATu�� ����6�r���@E�B���r/���56`l���dc?2�j?��X?(�<�x�>��������Z���A����@~��`������i|�5�GA�\�B�9<��KSAa{S�|�@k��@�*{�FǢ����տ���P?ROC22 i/H8�� m�%������z#�����@z>I5lﾓ��[�>�����)��A[��I�1@��@
����(�H��7"BGPOA��o°�C���SY�����x������C���P@S�״#?555>?G4� �� 2���o�?���?�**��c��>����>���'.�,^���:�A�
�@Ήc������R��v���L�B?y@�B��½:��CxXN�/���?�P>pK���?�7B�z��B��O/a!P1g N6O�
��3F���1@���@��$��.3�q���7�'.����n-$A��>(��A/V!B�[��A�BQA���B>��B����Cd������?�*?����? �`©Cf��O�Dh/�M�3E�>���?�V�?�zѿ��P�N����v^����;R�F>��ƠADm�B��O_r�A���B=���������Cd��n'.���?�6��=�O�>c-�K�.I�¥5�2�_�EO+��c/��%�mC�@?��4��?W�����@V|��V���
_&���f��A�h!@*����!?�$lW&�D>A	����V�����L�`bׯ���h��M�}A7�p��h`>��y�@���sjS1�05_DR_T2�0Ng �o��NT����3FI��?�����~��-���SAe�`����%��BP�@_<B�oA���QWr�}A��yA����=ϧ>��]ߟ���#n)#�wA������A�2@�+���W��sjPOUNCE_Se/�@�T�TI�%@��;���+���e�:?j�����
�'.��4P���'A5>��@�/��@'ݰ'.����o?HA�P��B�mS�Y�fíe�'���@(xf��!k�@h`�@p=�~�38PICK|p|�o�JT�Dg���/׭�jh��AJ�s@;&��(�P�&.��w��-�%�A��۸I@���?k�)W�"�A�:�?��3��Q���\n�9;+'.)�����5A�����V��@h���@�}!G~8o_PK_�N8
���T�E=3E;U?5�7W�#P���+���LA�����a�<@�p�@G�q@�"��W��B�,�����A��a�z�lo��6��#n��X����B������]��V�����ß՟�� )���n3E:z����:��l��P���԰WA��� ��z@�'<?�J�@\�TG�Y��_�Ec�g��kk�]P�2¼���B�&��S�4@����C�7������͢����< ���9�S���Q�( �d�h���A�k����@�2�?}O?�R��S��[������b}�g���6�5S��G~±��B��@�O5�@M�3��=x�]�ȧpVۡ���������jaA˒	��3� F�s@��￑�[��_�(�c�{?�]Pa.s�����B��w����0@�T+�C�BZ�K�d�Ǩ�Ӧ���m�^�=����<�5U���b<_��l�A�L�����@��@ss�@Q,^�ϑo�B,�������b��k����6����&���f>&��<��q` @�Y�@2�soa!/�	��+��E�3Eo�5��=���<��[������c����A8P���
�?�bo��9q���ߐ�B,�������b?�k���6�[�������?���H��@9�`@uz\/�����Ӧ����;:��>2�<�'�(�����\���K�hA�9�N�o� ?�����1?�j�S���&B,��������f	��l���6o�S�?��»B�?/����?0;Φ��M3����3E���m�M�\>�*��8�b��U湼�@��9�A��(����@WSQ�`�@/Ơ?�aRB�+���8��i���l���5y�m�!n�¶�VB�����M�A)���M��������F�Vx�`?9�/�(�=a��罍0=�F��@���A��<��(@�Q�=�D�@*�%U�+ N/ �3 �7 �Ǝ�6�E���B�D���R��A6�f�
ߜvZ��OC1<?��3Eὡ��>�\<�_�'_�!��B�A� �A�����^��@A�������Z	B�*W����r��g�|�k��7��;�g���O�B�����NR�Ac��@��67��./�4�3F�T?%W����=��b�e;�yd��A��A��V���(�@���Hbo�DP���X����w�g����k��7���>�����eB�v��\��wA]��@p���"K�@-���z���0^��J���=y����W~�� ;9�C�#n�VA�������AK?=�AR���m��&'J�E����C@�U�0���֕Jn��o��¿��B�T���|��O�=�ĚG~2Yr46�O¬������M����� �?dT>���e=� ����n�a�@��Iӿ�TA��4>BX
 @���c>%�*���-�����@�����7s���~��r���B��U�;��Q¯��K���G~4%��?�H'�T�������;�=�#>z�:;:T��9��ſ��� �����0��i߉����m�Y�R@�Al��a�����?����~���AQ��B(Iv�A���B�u�A�k��*Up9�YrCOMU~�(�T��D��<���G�3����C�%<�@������N;	�A��a�
��@���a@�c5?�����n3�B�(;[������b	2�i�v��4���Uf���^B�����e��.�@~�	,Tq6�32�/Ti+�T����vQ1��?�H���^�� �d��m��Af%��0���]qA�I�@�N�c@��	������rd�p�A�֧=�U��p���KC�=����*W�@��	�@�4A?���dµ�-��&Q����wRk�?�ٗ��Um�� ����[b�Af�K�������A�`@Ew�u@�������tk�p��`�=����p��oQ�5A���9Q=@{��@�xA���bh"��Q��{����������R��>>�R>��_)�n����h�`�7wQA�g[��.��9��B��C�q����K�Ba������ºS�������zm��UeO@l���sA�,��瞩I�/!C22� Io�{������!�$��l�);�;�Ӗ>)�H�������9A{� �;��	A���[��˯��L(s��w�P�{���ރ���M��}��*{����A���­��V����O׋}��s��~�9=&{�<��h�'B�=���=�
���}���Z�����A��@B;�|�����1���}B>�
�o���B0N�@����®�����G��h�A"���@�=\?��@? T�-7
PR�0PRMŏ�x���y���2�:=�P�V�>�b��g�w���t��������<Ac�9��!5�豟�����L)�o��B$��B�*��t�)x��Z��@��]@/��&?�/$@�?ґ@dQ�S�e��u_L� ��}�����A�;���\S��;�
ͼ'��.�`��������Ad�w��:R�@��3�?��,ׯE���p zB$�+B��3��0)u�U�ށ@�A
��!?y�?�!��@��@*�'�9��]��vS����i�A}P�>A��������A_�8��\�9/���_�����˞A�I�1��e?A�p���Be^��<=��B W�B���£[��ǽ�ܓ�w�A�����"A?�7�+�Bk���_50PIC�  }��J�wU6��'�Q�����U�۞� ��`S�A�J@�n��;�@5�/�����`�p@X���BW(|¶�ߚ�{8|�ޥ�����+�M�������?��@C]��!B�RIFICACA9O���wY���}�Ȑ;��u:009U�������ͨe����A���@ǁq����>@�&v�S�O�`�'@�Xq�o�sЍ��z=N�M��?�hZ?��?�T�v\a@�}!��߽�����f�\a��ш�����:��F9��\a��}=� ��7DA�֪�A�%����n�'�2�`���@hH'BW{'�s�v�{+�z�wA=����e���n?(`>a��<��n���yX����C�a@�@k�Aڰ��d��@�ފ�ە^�N�O���[C��2�AW����Af|s��iN��6�d�B%kA����W[�Ж2�N��A( �����nA����R=)BOަ����f�\g*T�{��?u�JI�� S���"l ��s��@���?X7�.�Έ�o��z�E�o"A.��c�W�AL��'�u@P�;��1B!��A�G�� J���~�$�^��[����U@|?>(`B��F��m�K�����@����A����kf@����۸�v�F�Ӵ��������AXl������Af�������������A��`���?A�N���Z�BL������Psm����@Uk�@D�����p���9�d�O����@A�>G>D�v�χX�h�f��S�H��AEt��<�f{���M��诮!����'�An&�G?jF�?h��?�K���/�0sm����^?�?��:�@����O�@� ��4A�'4� ࿞2�Ŀ��K/�i��?�/AA��<��k E����Y��������r	@��?#�H����>a���z���/��w�h�?z����S���|���~W�AfR������צIA�P@D�@;|��+ZZ�t]�A���A�ՠ�=���`��p0�/�0�?�����@p�@��vA?*;�`�4���fO�x�.?1��?�%��^����
�m_��AD݆~�ќ�����Atp@>� @�����@�?�l,A�$A����=��X�׿�\���3O��Y��$������q@*a�@S?&'�f��COUO�:_�y�5?v$��C?�l�\a�������m��ADТ�7������,pA�`@�|=@����}�J��O�O7���R@�^�����@O�g@��\`	_)_o��z;�?u<�X����{ٽs���<�s	�?��!�9C��μ���A����f>��Aan�@�	�^$��A�jB���������7�L����MO�5���ú�B������q*��z?�ŸBo:S10_7_PK_�N`�o )#`�?u����?��#����y<��A>W�[�<�"����yA�6~��U[cbb�:@
���oo��AjU�������_I�7�7�`%O��r�²L9B��h��-�� ��t���X�����zT������=���A>�[?�u�<�����8���B����(�A������?���@w7���A����FBM������:�C���z��A,6Ͽ#�����O������	�DRO�P�0�?�kT�c�X�X�9�;�\S�;��b!�Σ��@1����A�%r��,B�@籈��1�B����BM�U���17��C��J�#�5�2��_!���d0���-t�`�/��Տ�����>�4?0�S�>sQ�p�e��E�������ܵgAi��,�%:��@�^[C���R��I�ZA�5���$y���9�C����^@;��@ﳳ�?�ѕ��'v���Ъ��s���X����w�n_�>��R?2��>s�A�k�Ͽ�(~�����+��An���?�@Ơs@<p����\�I�A��=M�$lI���;�C���?���@�h>�O��xy� �~H������c����$�<��="���<O����н���O9q����>pAr!��;�3�@��J@Y��L���I���A�&��$��\��6�C����#.� AC��>�о�Ǣ�?<߿)y]�y��8N��������U�5�:빹�\�S�9R�p���=�u��{޼�����A��c�؀@)���@z{g�
���I��A����W$�釰[���O�R�?w�������X�,@���9�b���ɵ�ozU	�v���n>RZ-=����>
܅��?���#7k����OA|��߂�Ơ@S�X�����K�A��V��)ء��̒o���OE���@�oW@��/�8�Ϳ��?I�t�OMU�����`�vԙ+?�p�>��=�l�����E����O����q�AB��J$l@�:@�{\�Z˓/I�8�EA���"��2��+�C���l?���@Č�x@%3�=�aM��>���w� x���̌�5��5����l���2���IP��8(�<��N>�����N�c�}�@ތP�g]q�]�%��n�2����z4@Ǔ�)�	�ס�O����9�B��rfA�:�����B ���{7TY3�Ͻ}���0�1��H�=;^�/�9� :8� G>���v����A�O⮽`0� ??�C#%�@�����%x���W��p��k��O����S�MA�����O@��5����R�n5_DR_T�2�o 
OT}M�o���������:�>󼮵�ݾ�<2#��Aj��+A����7�?A� A��n��E�u��$���9�������AɈ�&�����@Q�������\�B�������7����?�"��n2���41п�}d��5>���?`��N�x��=�\��>Tqڼ�K��Nl2�A`���?��AP�Aϻ���@ _���9�i���[�Aʞ�&���� s����²�SB��T�֗O:�<@@\�|71K��,}�6��);M�5A���o|8Bu�O�Ǝ��2[���Cw߭q�f�����������<�n�<_�{�4�j�AI��,A�A-�.��A�}AT?��?����$���:<��M �Ar��'t���2�Ҵ?�£�pB���������˔�@����c/}/�s��5`�=�|�=������G���<�ӗn�\�@۸I�����AUYA���r��/ ���;���-|A��g�'����8���P=o��+@Ԡ@:[(@� �����+?�1�8N8��uo��]����!���SＰ[��A��<R4:��R.hA�z!����A\цA�i����On �:d�*��kEA���&�H��9��s^P��t���A��?�`� >�����ɀ�?�q O(N���SV#�m?�����\�ž�mb��m�AD���s^����NS�A��@v��@�V!�~7D�_�^[�_�P�\�@�ǲ�'Y+�@T�v@�1��\���_�VF?i�dZC���ay���羒�q�=�~G��p���aFn@������A�Ʋ���d@�f�@��W]�	�u�D=�`���n�k��S}B#�bο�T��x���x��?c-K�S&'�E�l8?�o��u}�f�����`�S�=\��տ�A��U��R��Z��(�A3��ٿ�boA��&CQW]Bf`��f��BVvG�A0��!X�C:Ƈ>|�����?�l���x�h���g��?3�ɿr 'Tw~Q�f��կ��o2`�ﻁA���^>�����bA�4�V�b[�7�Q5�of_%�@����+�?����������y�mK
�Oy�6�Oz|��6��{�쁑��?,�~v+���$8@��@�)������:����A�a�3�����m��׋�6�:A������Q��T��R�߰��>5�������A$�����/$@c���O�07_PQK����"[��_��`�7#.>�[��=b\���ߏ���c����#x�Aj8�����>@Oj�a@Ч�L�A�����\p���v�NɎ�8'��b0�����"A{����-K@��L�>���韬f���_���l�<������� �����>3'=3�.@&������A��@:R���&�����{�F�A�{���/���F���O�6^����@������AL[������@
Vʿ،ڰ��	�¯-��_���#=L=��:��D��U�?�Y�>��@]�zE����A�J�@>���T ���O�A�A��c���'<���)n�P������e����hZ?�m`�!{������⟯豯��բۦ(#z�=��(�JT��h�i?��>�8��>Z���z@1\���P���
��#�>��A�H����m��ʅ<�Q7���w�@�?���?��>v��?.m�S״s�腿j�բۦ,s(�=���x�e��?��#>��禎@^[C���A�+�@H ���w��*����;VA�3����r$��پ�Q�n�O����Y?�� ?�֌��*a�??�� ZJS��l�Ϩ_�9L�>���s�O
����f?Kr=��Y�oa��QA��:�@���d�7������>KA�������������Q��ב�_W]����տeARB��D��H��:�I �4ߦl�_�K�>��$�W)����:?K��=��yxc��q�M{A���*@G�q�p��`���>QA�dP������ɫ	�R�m���Sn9�����hA.�R7�?�7@u?�ڿ�.��ߕ��_�"3�>�Y��D��ނ>�?U2=ҌK�p���8A�/�@oK�h�<�	��N��TA�.N������}7�R����G��!�����T�AA����@}ɿ�Y��ט�Q�
��3ۦpٿ�\���C��`�s?7C>����>i�,����A�Q�@�WSQ��0�1��G�3�A���������� [��SG0�W�Sn�@��W�P�@rp�?��=?t`��X�-��բ@۩�\�Y߿U�����>!�!�>-#���#:A���D@Cz�T��W���h.<�A�(��������#��S���n�������N?AD�L��M�@s���)y]k}bբ�Rۦv"���ſ׬ɾ^�e?2�>�`��Ͽ�"��A����@R\���lk����'��A�]��;���*k�T>�.��~T��JA6�3���ϧ���L1/Ч�Uۦ�4q�"x�t� �޾E_�l?U��>��k�>n-$���A罺e�Ҽ���!�A�������2��<��T�UQ�~�����7|A=V����P�"i��/%/
?բc_���ΌA���#��5��
�>��Y�=��@�C�x���A����g�Ew��8��/�A��r���&����6�U	�b����r�����_A;�1�3�ґ�2C��/�/�?բg+��:&{���!߹R�p9�`�d�A?[���A�ҿ�?�����`��h0k? A������X����a�T���Z��T @D�x�@�g����<������Ġ���B�0i�j��?�u>�ҟA�b�O:����#A`���?Hbo�D��v�=�v�O@�A�Ƿ��}H���o_@��YF�wA����A���
��m�@?�QB@*ʟ �����Ol+�ȫ=���W���Y��}<�q&�rA�g��?��R�~��O@A�Ԕ������?_@��7P�������A�Q�ſ��@?�;?�B�Z�ٴg�^o+麝@����P�:�=:�+N�_�pY��A�W�>o"��VrS���L��_�Q�!��^C/���_@�7Pv���B���AI����Ι1?ŸBL7oݒ46Po�]�3��<Dps�C���@�p�_�T�",A���c>��ٿAZ}�����o� A�����K����_@v�7PHo1ÿV����v?�=�3�&ݒ13�?�]��W�?��?����9@:`�ӌ��Ш��A`����1�P�L�� �A�+��G���/_@57P�����҄7E~�1@�hD?a���ԏ#����q�?�D6��a7������v���6A\��G�Q7A�Pc� �A�.���B�M��7_@��X�NTdU?A��c����<�=ؗCOMU������E��m�	���
qͺ��:T;�+:����o.���I��,A�h�@?����fD3�$�Y�7��A���_��!��ħ���U�g��o-�b0��f�>&A_!��8��@�<߽�}��?y��7�Ö��m����f���q����F:���ߟ�0�"�"���
?۸I��Bϧ��2�J��A�^�����'�_%�U0/��o.���0��u���?��?���7��p�[�m�R��2���E������!���8���@�p�����|ε��=�_EA�`/��� �@�`߮#A����Z=�h��(�y�/�zzo.P��P�?��>�Ǣ?
V�?�ܤ�����Ƨ]p��p�ǿ�����Q??]��F�o.,B��� HA��A@'�ݰ�� @�����#A���^PJ�iWp¿�l��/�^�?�1����9�A�E��?FǢ�?�NX@i����)��ԧN��]���������?L���7_o.<���A����޴`@X����A
��W����hA�8��.�ߓ>�h�����ADO���1?��P@X���������%�٧Q���c�c����6���?N?3�8�Qo.�p��cA����@Q,^�a�<�@A�.Ck�A$��Qo��f�+#_��-�շ������!�҆��@.���ߠ����Sr�o�ftٿ�}����{�?O��9�o. ����A������c�9@��/�	�A71��J݈�e}~���9�,�t�o��@�8���<�-�K?�E�@<M����v����R��Ŀg�X���E`�Čt?M����:Do.7�����VA��ۂ@�`�p��@.�*��BA�O��D9w��d&�����+���>�Y�����AJ6i����@+���qUC�Km�n��K��@7�Z�@'���5��@?=(�����5�AYN?�{Β�a>��>����A �b�F���d�j���,H�.b�XA�{���O_@T�#����,'e��2+��$SERV_MA_IL  �M��Pp7OUTP�UTBP@>7RV 2Is&S_�  (�DKPpI73PpPp�A;$�7SAV��e�TOP10 2J�� d �@b �!�@�Pp-6 u%Pp
�B ~ }SR6 &Pp��@R 2  ��� sPp~# *RPp1 .! .O"�E r/$�O" -'O#�O$� 
�A[ eR۹�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O��Oݳ�YP��F�LT_CURGR�PBPpM=TI�DX  �M ��#|_�W:WNUM�GWL
:TDISF�UFP�1]ERR"PB!n~!9U�PTI�W�sS`:TON  k_=oKj~:TSCH 2K۵=�R
�o C�MQ��Lt�o�n �U�o�o�i�o; &_J�n��� ����%��I�4� �R]�p�{o�o�ȍ�o ���9�&��6�\�G� ��k�����ȟ���ן �"��F�1�j�w�y� ���������ߏ�� U�B�-�R�x�c����� �����Ͽ���>� )�b�Mφϓ��Ϩϳ� ůׯ���(�:�q�^� I�nߔ�߸ߣ�����  ���$��!�Z�E�~� i��ϱ���������  ��D�V���z�e��� ������������ @+=va��� ���������<3� `r������ ��/�8/#/\/G/ Y/�/}/�/�/�/��/ �/+X?O|?�? �/�?�?�?�?�?O�? 0OOTO?OxOcOuO�O �O�O�O�O?__#? 5?G?t_k?�_�_�O�_ �_�_o�_(ooLo7o po[o�oo�o�o�o�o �o_!4?_Q_c_ ��_���o���  ��D�/�h�S���w� �������я
���.� ;=�P�[m��� П�����<�'� `�K���o�����̯�� ɯ��&��J�W�Y��l��$SFLT_�WAILIM  �l��_�  蓷T�����REC_GRP 2L����wʐ x?���;�)��Mχ�ZN_CFG M�Aϲ����l�ݲN���ɐ,B   A���l�D;� B����  B4l��RB21��GTDSCH 3O���� �   ����%�7�I��x�]߃ߕߧ߹�x����k� �6���{����HELLr��P��l�F� ��o�l�%RSR v�w���������
� ��.��+�d�O���s�@����������Ǒ���"Ǒ%��"l������_�t�<^_ )�l�
2t�d����|��)�HK 1Q�� �>���� /*
c^p�� ����� //;/���)�OMM R�7�w/V"FTOV_7ENB�� ̵��OW_REG_U�I�/��IMIOFWDLb Sf.���"Ļ��"�	�'��OU�T����<�����+?VAL ?�#_�UNIT�#b6̹L}C-�IO 2T���y/�?�?�?�? 5/O0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�ˏ_ �_�_�_�_ oo$o6o�HoZolo~o�o���2SoU 2U�<\�� �t�q��b�e�o��o>ǿ�  -?{) _M�qvO��������gLERR� 2V��� � �J�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ����\�n� TRY�'�%��1MISs�2W�< ��{O�χȨ�QqE�8�` wr����x������7�� �_IRD_MA/P  ������)�MB_HDDNw 2X� � �e�ݡ߳������߀���7�C�o��O�N_ALIAS {?e1�( he�o ������������,� >�P���t��������� g�����(��L ^p��?��� ���$6HZ ~����q�� / /2/�V/h/z/�/ �/I/�/�/�/�/�/? .?@?R?d??�?�?�? �?�?{?�?OO*O<O �?`OrO�O�OAO�O�O �O�O_�O&_8_J_\_ n__�_�_�_�_�_�_ �_o"o4oFo�_jo|o �o�oKo�o�o�o�o �o0BTfx#� �������,� >��O�t�������U� Ώ�������:�L� ^�p���-�����ʟܟ ��$�6�H��l� ~�������_�د��� � �˯D�V�h�z��� 7���¿Կ濑���� .�@�R���vψϚϬ� ��i�������*��� N�`�r߄ߖ�Aߺ��� ���ߛ��&�8�J�\��������m���$SMON_DE�FPRO ������� *SYST�EM*u�8��R�ECALL ?}~�� ( �}z�@A�S�e�w����� /� ����������> Pbt��+�� ���:L^ p��'����  //�6/H/Z/l/~/ �/#/�/�/�/�/�/? �/2?D?V?h?z?�?? �?�?�?�?�?
OO�? @OROdOvO�O�O-O�O �O�O�O__�O<_N_ `_r_�_�_)_�_�_�_ �_oo�_8oJo\ono �o�o%o�o�o�o�o�o �o4FXj|� !������� �B�T�f�x�����/� ��ҏ�������>� P�b�t�����+���Ο �������:�L�^� p�����'���ʯܯ�  ����6�H�Z�l�~� ��#���ƿؿ���� ��2�D�V�h�zό�� ����������
�߯� @�R�d�v߈ߚ�-߾� ���������<�N� `�r���)������ ������8�J�\�n� ����%����������� ��4FXj|� !������ BTfx��/ ����//�>/ P/b/t/�/�/+/�/�/��/�/??�#�$S�NPX_ASG �2Y���<1��  0b�!%�/c?� ?�-6�PARAM Z�<5F1 �	*R;P�$� �(�4��/0OFT_K�B_CFG  ��#B5,3OPIN_�SIM  <;��2OO1O;C/0P�OTTSKINF�O 1[<; g=R8~O�O�O�O�O �O�O�O_ _2_D_V_�h_z_�_�_�_�U/0R�VQSTP_DS�B�>�2�_$;SR� \<9 � �& STYLE�108_TC_R�02  04 K�U�5�6)6TOP�_ON_ERR � Qf�8caPTN� <5�`�A_bRING_�PRMmo /0V�CNT_GP 2q]<5�1H1x 	�_��o� �o;(7V}D�`RP 1^�9�0,q8Av�� �������*� <�N�`�r��������� ̏ޏ����&�8�J� q�n���������ȟڟ ����7�4�F�X�j� |�������į֯���� ��0�B�T�f�x��� ��ÿ��ҿ����� ,�>�P�bωφϘϪ� ����������(�O� L�^�p߂ߔߦ߸��� ������$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@gdv�� �����-* <N`r���� ���//&/8/J/�TrPRG_COUNT�6�a�5v"'ENB�oq%M�#�4��/_UPD 1_>kT  
_/�2 �/????:?L?^?�? �?�?�?�?�?�?�?O O$O6O_OZOlO~O�O �O�O�O�O�O�O_7_ 2_D_V__z_�_�_�_ �_�_�_o
oo.oWo Rodovo�o�o�o�o�o �o�o/*<Nw r������� ��&�O�J�\�n��� ������ߏڏ���'� "�4�F�o�j�|����� ��ğ֟������G��B�T�f�������h,_INFO 1`�%o�  �] �����'��<����-�8�CL7�A�#�Ay�u�<�fG���ￎ��g,YSDOEBUG� � ��d�)��SP_PA�SS�%B?��L_OG aݦ�#���鱄^�ܜ����  ��!��?UD1:\ϴî�в_MPCտ P��\���2#�~5�SAV bؽ����X��SV���TEM_TIM�E 1cط� � 0 �+���a%�����������#T1S�VGUNS� �%'��%�6�ASK_?OPTION� �%t�!�!V�_DI����/r�BCCFG #e�)rҭ��X���`��4����� A�,�e�P��t��� ��������+��O� :�s�^���������������� 9K�� 6e7��%�� ��(���%Ll� Pvd���� ����/</*/`/ N/�/r/�/�/�/�/�/ ?�/&??J?8?Z?\? n?�?�8u �?�?�?�? O�?0OO@OfOTO�O �O�O|O�O�O�O�O_ _*_,_>_t_b_�_�_ �_�_�_�_�_oo:o (o^oLo�opo�o�o�o �o�o �?*HZ l�o�~���� ���2� �V�D�z� h�������ԏ��� �
�@�.�P�v�d��� �������П���� <�*�`�x������� ̯J��ޯ �&��J� \�n�<���������ڿ ȿ����4�"�X�F� |�jϠώϰ������� ����B�0�R�T�f� �ߊ���v������� ,��P�>�`��t�� �����������:� (�J�L�^��������� ���� ��6$Z H~l����� �� ��8Jhz �
�����
/ /./�R/@/v/d/�/ �/�/�/�/�/�/?? <?*?`?N?p?�?�?�? �?�?�?O�?OO&O \OJO�O6�O�O�O�O �OjO_�O _F_4_j_ |_�_\_�_�_�_�_�_ �_
oooToBoxofo �o�o�o�o�o�o�o >,bPrt� ����O�
�(�:� L��p�^�������ʏ�����$TBCS�G_GRP 2f���� � �� 
 ?�  �%��I�3��U�l�~�g������şם��h��d����?�	� HC� ז&�ff$��ו�A�x�A�N�D)�ז���l�ؔ`�B4N�P�b�Ln���-���y���ޭCj�����333וB�Cޯ��י�i��4�ؔ>�v�X�B�n���@-���-�ܵ� ��̿�7���b����dȰ��	V3�.00��	rc;2l��	*�������Ϙ�G�?��33�X��d� 8����  =�\��Q�Z��JCFG j����Z�+��&�Z߯�������ڽ��� 	���-��Q�<�u�`� ������������ �;�&�K�q�\����� ������������7 "[F��%�� ��j��) M8q\���� ���/�#/I/� ԏn/��~/�/�/�/�/ �/�/?�/4?"?D?j? X?�?|?�?�?�?�?�? �?�?0OOTOBOxOfO �O�O�O�O�O�O�O_ ,_"�D_V_ _v_�_�_ �_�_�_�_o�_o:o Lo^oonopo�o�o�o �o�o �o6$Z Hjl~���� �� ��0�V�D�z� h�������ҏԏ� �
�@�.�d�R���v� ����h_֟�����*� �:�<�N���r����� ̯ޯ����&��J� 8�Z�������^���ڿ ȿ���"��F�4�V� X�jϠώ��ϲ����� ����B�0�f�Tߊ� x߮ߜ߾�������� ,��P�b��z��J� H����������&� (�:�p�����R����� ������$6H lZ�~���� ��2 BDV �z������ /.//R/@/v/d/�/ �/�/�/�/�/n�?? 0?�/`?N?p?�?�?�? �?�?�?OO&O8O�? \OJO�OnO�O�O�O�O �O�O_�O4_"_X_F_ |_j_�_�_�_�_�_�_ �_oo.o0oBoxofo �o�o�o�o�o�o�o >,bP��B? ��H?~��(�� L�:�\���p�����ʏ ���� ��$��H�Z� l�~�8���������Ɵ ��� ��D�2�h�V� x�����¯���ԯ
� ����.�d�R���v� ����п������*� ��T�f��>τϖ� �Ϻ�������8�J� \�n�,ߒ߀ߢߤ߶� �����"���F�4�j� X��|�������� ���0��T�B�d��� x������������� P>tb�� ��x���
�: (^Lnp��� �� //�6/$/Z/8H/~/h.  � �#� �&�/�"�$�TBJOP_GR�P 2kp%��  ?�Ҩ&	�"�#m�,��x  ��� �,^�% ��� � �s � ��$ �@� �"	 �C�� X6Qp�D����%�!t2&f�f|2q5}?�6<9�]X1?��?L��Ͱ1BH  A��n7�?�7D)�\�5d2�Sl>Y�0�A�1	O �2�0>̿��<���1?�333?f�0A@B�  B �?cO�?D5ml>-D�6�M8�1�1�1Af�<B�E�� CQ@LATO�OCj��V�?�KAA)_;Z�;ć�B�@FQ��@�O�__�_�H�_�^<��\Z���l_o�_�_ t6u44AHoN0EAE@4B�z�J\R�T>���C4N@�o�oBo �I�o�o�o�o�o- LfP���� ������M� f凨&�p�t5	V�3.00�#rc2l�$*���$�!����� F� � F�  GX� G7� GR�� Gr0 G��� G�@ G��� G�\ G��� G�` G��� H
� Hd� H" H.�� H;� HH2� HU�ÂE��� È �F@ �F�Fj` F�?� F� Ȃ���� G$ G��GV�ۃ�� �G�L G�� �G�h G�� �=u=+8�X���z�/����zg��?�  L5�@��.CPPACT�SW  �)��IoR np%�!�  C�0 �SP�EED o*� �;�]�  }�
���_CFG p*��!��$�l� �_CUR_ID����6���EXT_?ENB  ��Х���HIST_B�U 2q�+d o}��j���������j�fr�Uj�j�j�j�TQDp�&j�,j�2j�U8j�>j�Dj�Jj�UPj�Vj�\j�bj��hj�nj��3�"�3�(3�.3ȍ`5�:�3�L16�F3�L3�R�3ȃ�6�+5:�d3�j*3�p3�v3�|3��P�5�k6;��3Ȕ3Ț�3��D9¦3Ȭ3Ȳ�3ȸ3Ⱦ3��3�ʪ3��3��3��3��*3��3��3��3�̀!�i�����&��*&���$���(%���$�6�<�堨!�[��N�T�Z��`�f���%�r��x�~��������������������f����Ր!�������������_MAOX_AN��Ǯȸ��SPD��rȭ� �^��:�o�%��8!���NUM��!�̩
��OUT 2s�+
 �����	�� ������ *[Nr��� �ZERO����%?ESTPAR;`��7�� HR�AB_LE 1t�+��F2h������*D�!�	�u�| � �.�r�| �`N"RDI/��./@@/R/d/v/�%�$O�/�
;?&?8?J?\>"S$�/��@2��"�N�"A��0��A��0Z�BA��0�1A.���BA��0�1A2��2A��0����0�)��O�O�O�O� �8���A!8��!AJ�	r�A#8��!AN�`_0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�oC�0�? (,��?�?�?�?�/�/��/�/�/�""r[ U*��p@_ ` "��u*�u��� �IMEBF_�TT��u�H�VEЪ�`��[�E�R {1v�� 82�ro " ?�  ��7�]Pm (�����ҏ��� ������/�A�S�e� w���������џ�,� ��b�=�O�a�s���F�� ����ϯ������ �̖� �2�➪��d�v� :CG��������Կ���
�ϋp2�D�V� ��l�~�����P���Zw�@����?MI_CHA��U� �� �DBGL�VLQ��ET�HERAD ?j�u��ip0~��:e��4:3b:�57:e6 ~�7(�ϋp��9\�R| o�!��!����H	~"�SNMASKj����{�255.�0�f�.�@�R�d���O�OLOFS_DI���%ORQCT�RL w��Rsiz��qT������ *�<�N�`�r������� ��������$���G6k�PDRA�M%�x��d�s��o����  $6HZl{  ��)������E?_DETAIHؕ��PGL_CONF�IG ~�����/cell/�$CID$/grp1{/+/=/O/a/ +ħߌ/�/�/�/�/�/ u/
??.?@?R?d?�/ �?�?�?�?�?�?q?�? O*O<ONO`OrOO�O �O�O�O�O�OO_&_ 8_J_\_n_�O_�_�_ �_�_�_�_>~}�_4o FoXojo|o�o�q\�o�m��_�o�o!3 E�_i{���� R����/�A�S� �w���������я`� ����+�=�O�ޏs� ��������͟ߟn�� �'�9�K�]�쟁��� ����ɯۯj����#� 5�G�Y�k��������� ſ׿�x���1�C� U�g����ϝϯ������������Us�er View �)}}1234567890(�:�L��^�p߂ߊ� ��+��C�.�D��@;��B����ów���2 ه������"�4�F� ��^���3�ߔ��������M��q�4 ��H�Z�l�~��������q�57��� 2 DV��wq�6��� ����
i+q�7�dv�����q�8S/*/</�N/`/r/��/�" �lCamera�/�/�/�/? ?2?bE�/\?n?�> &ߚ?�?�?�?�?�?��  �&���/DOVOhO zO�O�OE?�O�O�O1O�
__._@_R_d_�/� �&���O�_�_�_�_�_ 
o�O.o@oRo�_vo�o �o�o�o�ow_�W6�go .@Rdvo� ��	����*� <��o�WK������� ��ҏ䏋��,�w� P�b�t�������Q��% �	?�����*�<�N� ��r�����៺�̯ޯ ������WR��`� r���������a�޿� �M�&�8�J�\�nπ� '��W)�������� �&�ͿJ�\�n߹ϒ߀�߶������ߓϥ�9 x�-�?�Q�c�u��.� �����v�����)�P;�M�_��	�%0�� �������������� *<��`r��� �a�s�� �+^% 7I[m���  ���/!/3/� �%'K�/�/�/�/�/ �/��/?!?l/E?W? i?{?�?�?F/���[6? �?�?O!O3OEO�/iO {O�O�?�O�O�O�O�O _�?�5�k�OW_i_{_ �_�_�_XO�_�_�_D_ o/oAoSoeowo_�5 k�o�o�o�o�o �_ASe�o��� ����o�5כz/� A�S�e�w���0���� я�����+�=�O��}  �y~��� ����Ɵ؟���� ��2�D�   �qD�2$D�^V?��v�@�X�B�s^��q��?�CD���5���@Jo�B0�P�DЖT�?���B8P��n�����=m��C��B�H��T�@�x�����+�C�.�D��@F�B����ówĪ�B����D�y�?�
�Z�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲�����p
�p(  }�r�( 	 �� ���� ��D�2�h�V� x�z���������
�:ܪT� ̞�O� a�s�揗��������� ���s>�-?��c u������ L);M_q� �����// %/7/I/��/�/�/ ��/�/�/�/?!?h/ E?W?i?�/�?�?�?�? �?�?.?OO/Ov?SO eOwO�O�O�O�?O�O �O_NO+_=_O_a_s_ �_�O�_�_�__�_o o'o9oKo�_oo�o�o �_�o�o�o�o�oXo joGYk�o��� ���0��1�x U�g�y��������ӏ ���>��-�?�Q�c� u���Ώ����ϟ�� ��)�;�M���q��� ��ܟ��˯ݯ��� Z�7�I�[��������ൿǿٿ � �@  ����,���������+frh:\�tpgl\rob�ots\r200�0icf�_125lif.xml� �Ϥ϶����������"�4�$���>�c�u� �ߙ߽߫�������� �)�@�:�_�q��� �����������%� <�6�[�m�������� ��������!8�2 Wi{����� ��4.Se w������� //0*/O/a/s/�/ �/�/�/�/�/�/?? ,/&?K?]?o?�?�?�? �?�?�?�?�?O#NEȝ{� �P�8?8�?�#KbO #O^O�O�O�O�O�O�O �O_ _"_L_6_X_�_�l_�_�_�_�_�_k��$TPGL_OUTPUT �.��.� F@�DߑC����Q@'�A���C�w�*�ē�vDZ�D���`@��B�?  õ>.ewo �o�o�o�o�o�o�o +=Oas��@�����wF@��P�2345678901��*�<�N�`��h�$��Pnosel�ect**�*�)�9`D3VS�*���a9`  |vH�Bzk5?���+��D�EB��z��*��1������ hh0B���$��*��܀�.B������%� 7�I�[�m���r����� ��П�z���}��� /�A�S�e�������� ��ѯ������+�=� O�a�s��������Ϳ ߿񿉿��'�9�K�]� oρ�ϏϷ������� �ϗ��5�G�Y�k�}� �'߳���������� ���C�U�g�y��#� ����������	���� ?�Q�c�u�����1���@�������}AA�GYk}���@�HO��NJ ( 	 �A/ eS�w���� �/�+//O/=/_/ �/s/�/�/�/�/�/�/�???K?9?o?�v� D@]Bw?�?�=�?�?�? �?O!O�r�?JO\O�? �O�OpO�O�O2O�O�O �O_4__$_j_|_�O �_�_T_�_�_�_oo �_*oTo�_Do�o�ozo �o�o<o�o�o,> bt�o`��^ ����(��L�^�  �����r���ʏ4�F�  ����6�H�&�l�~� 菢���V�ğ�ȟ��  �����V�h�
����� |�¯ԯ>��
���� @��0�v���򯬿�� `����ҿ�*ϔ�6� `��PϖϨφ����� H��߶�8�J�(�n� ����l߶���j��������"�4�:��$TP�OFF_LIM ��0� �1���O�N_SVS� � �e�P_M�ON ��5�g�� � 2�O�S�TRTCHK Ƀ�5e�Dm�VT?COMPATz���i�VWVAR 儚�'�~� R�� ?�� ��O��_DEFPROG� %��%ST�YLE108_T�C_R0����r�ISPLAYZ���o��INST_MSK�  �� ��I�NUSER���L�CK��QUIC�KMEN'��SC�REF �5�tpsc��a hf	e�w _{	ST���e�RACE_CF�G ���'��O�	H�
?��H_NL 2���c0�.� T�,>P�bt����IT�EM 2� ��%$12345�67890�� � =<�///7# G !=/E+Q�/ �/H���//�/�/E/ �/i/{/D?�/_?�/o? �????/?I?S?�? w?#OIO[O�?O�?�? O�O+O�O�O_sO_ �O�O�O?_�_�O�_�_ '_�_K_]_&o�_Ao�_ eowo�_�o�_Qo�o5o �oYo+=�oI�o �o�oc���U �y��!�9���� ��	���-�?��c�#� ��G�Y���o��󏼟 �ן;��������� ����˟E����ӯ 7���[�m������O� u���믓��!�3��� �i�)�;ϟ�G�ÿտ �����������S�� w���R߭�m���}ߣ� �����=�O�a��߅� 1�W�i��ߍ����� ���K�����)��� �����������5����Y�k�4�S��|�9
�  ��9
 ����
 �����h
UoD1:\���K�R_GRP 1���� 	 @ ?Q;q_�����������//</'%?�  W/i+S/�/w/�/�/ �/�/�/�/�/+??O?�=?s?a?�?�?�?�?	��?�?ISCBw 2�U B/ ?OQOcOuO�O�O�O�O��O?V_CONF�IG �U�� P�./9_�GO�UTPUT �<U	$P��?_�_ �_�_�_�_�_�_oo�%o7oIo[oqPRe�gular Option`o�o�o�o �o�o�o $6HZ���p_���� �����'�9�K� ]�ldu��������Џ ����*�<�N�`� q���������̟ޟ� ��&�8�J�\�m��� ������ȯگ���� "�4�F�X�i�{����� ��Ŀֿ�����0� B�T�f�w��ϜϮ��� ��������,�>�P� b�sφߘߪ߼����� ����(�:�L�^�o� �ߔ��������� � �$�6�H�Z�l� Ua _m_���������� ,>Pbt�y� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/��/�/�/ �/�/? ?2?D?V?h? z?�?�/�?�?�?�?�? 
OO.O@OROdOvO�O �?�O�O�O�O�O__ *_<_N_`_r_�_�_�O �_�_�_�_oo&o8o Jo\ono�o�o�_�o�o �o�o�o"4FX j|��o���� ���0�B�T�f�x� �������ҏ���� �,�>�P�b�t�����>{������ʟ𴑣�����  Re�gular Op�tion R79�8 : DRAM� File Storage��K�]� o���������ɯۯ� ���"�4�G�Y�k�}� ������ſ׿����� �1�C�U�g�yϋϝ� ������������-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��������� ����%�7�I�[�m� ��������������� �!3EWi{� ������ /ASew��� ����/+/=/ O/a/s/�/�/�/�/�/ �/�/?/'?9?K?]? o?�?�?�?�?�?�?�?��?O�$TX_S�CREEN 1��̕����}ProdHo?me.stmObO�tO�O�O�O�	P�ROD HOME�N}��O�O__(_:_L_�O�O�_�_�_ �_�_�_T_ox_%o7o�Io[omoo�_mh�ttp://19�2.168.1.54�o�o�o�o�oATI TC! o^p�����o A� ��$�6�H�� Y��������Ə؏� a����2�D�V�h�z������/wizinstMOڟ�����"��HWiza�rd Top M�enuJUALR�M_MSG ?�2I� �  �INVALID �ARGUMENT� RECEIVE�D2|�DEC�ISION CO�D�GWAIT�ING FOR �MAINTENA�NC�ETip� Dresser� 1 Disco�nnect Of�f��ܫJamm�ed7ڨ G1 CurrentG�_o Lowؠܠ�d�(s) No�t in Aut�oէ �1 Mot�orI�Start��Z�l�oppv��STEPPER �NO��SET:�Watersa�v�Unable~G� Reset���2ȿܫPha�se4�ss0T_�4z�J�Acnow�ledged WSC1x�%�2ح2鯢��2	����2(�OBz�2f�x��˓�R���2	˗�����WT�R 1: WAT.��OFF0�2A�1�Mؠ|�&�Dum}pD�dvanc��SMz���Retracu�����y��ٯ���3�� T�������4���E�/��7�WN٬�k�L��3T	��3(�`z�3��(x����_��3	�۪0E�k�]���CS��4(�z�4�x���ꓳD��4I� Check <�F�PinF�����%Equaliz堯Faulװ 7�x|��)�High1�ؠCap C�hange ERWROR,�1�l�M��P�� Co�u.�� �Find���2�D�4?S�3��
�P�-���Search �Sens��ICoSE� ofb�^IOñTr�°lHy Anti� Cras�TM�_iRVisҲrv�鴤����3END/9.p://^/4RT1z/ 9 �/m/�/�/�/u�Key Swiqt`��N�UTOV��- iGun?/Backu��J�9P-@D>�z�H���7zoff �detq��* CH�| s nK�tohe c��ri0��  $z9�|�1r�emo� /őal�.�5 2 Ad/apt.ұi�0��� kN i�1��TD Verification�9� >�8samew as�1ach��� CZ?j8 ��ڠP@ogram� ��DISP_S�EQ Error3 ':Ol91zOj9�%yOk:7y�j9N �g�Oj9{��Oj9�4_j9>:_j8
�Z_j8{Pz_�_�_&���v�_j8y�_j:�# �_�)oj9��9�:oj8�>
Zo�_L�oj5��oj:*�o�j8o.�o+��omXEɔj9j9<1�	Z,o�p8�j7q��Yo,Z]��j8H�4.�j:�j8[�x;�j8-�[z�����U�Y_�o��2j5x�j:'"�Od\�j6ُk:z�8̊�j9�J}��MY*sڟL���A��_e��LTZ��+z�m�a"��K�ܯj5M>���*�M��j8G'"d��)t�Oj9����&j9ٯ˪幯j9g ��j8�?y��j9	���j8��9�j8AD:�j8g��Z�MYp�z��)
ƚ�j8_ �̺�j8Ko���j^f���j8���j8s��:�j8��Z�Nj8OBLz��	/y��j9��R��j8���Y?j9PN���j8�s���j8��^:�Nj8���Z�m����rj9�8Oj:����j8¯���j8�E9��j8����j8'SHE:�L�TY�j9'UG z��)S�j9�DU���*EY�j9�9��j9I���9���j9/�(Zj8'��z̩Nyo��SK:intSh;op?R8��8�O]?��8�?���8NU�:�8Ds_PZ�8X(UzΊ8=&��8�_���	IG��8Ts�#��8�)/f�8��)ɯY��)&��z/�8�59̚/�8H�2�/�8�����/�8�y���/�84?�8����:?�8;D<��$UALRMn@V�  ���1�� � 7 &�2�4�;p�7�7�?�2&&�?��?
OO.O@OOKz0E�CFG ��5c�0�r��@�U���A   B�ra_ 
 �p�xD��qA!(�T����O �T��]L�N ���@��O�w}T��r�O"�&T�Z��O$��T�\s_6aT��+P�M(/�T��{�D_/#T�|�i\_*pP�aAG�RP 2�kK �0�B�q	 @+�<5?�Y>���o9ȕ������6k�$�UI_BBL_N�OTE �kJT��l���5�w@�RDEFPR�OG ?%�; �(%	PRT41�PICK  20�4_MKZ�  �%S103_PK_T13N5�P eoPb��oyo�o�o�o �o�o�o0T�W�INUSER  �mZ^_ME�NHIST 1��kI  ( �(`��'/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,33,1 3a�p7`�r�	��-�?�� ��,�74�qR0�9 2 �������M�_���w7�rUNC�q2�,8Ǐ �2�D�ӄ(�ۏ�93{�ROP}1�p7 ,82K������ɟԃ._��e�dit�r.`50_���4��(�:�L�ӏ,i��t18�qO���33S�����ѯX�r���6�q4`�����2��D�V������38,2�������ÿտ� a�qE��/�A�S� e�`����ϡϳ����� ��x���1�C�U�g� �ϋߝ߯�������t� ���-�?�Q�c�u�� ������������ )�;�M�_�q� ���� ���������%7 I[m����� ����3EW i{����� �//�A/S/e/w/ �/�/*/�/�/�/�/? ?�/=?O?a?s?�?�? �?8?�?�?�?OO'O KO]OoO�O�O�O�O �?�O�O�O_#_5_�O Y_k_}_�_�_�_B_�_ �_�_oo1oCo�_go yo�o�o�o�oPo�o�o 	-?�ocu� ����^��� )�;�M�8O������� ��ˏݏ���%�7� I�[���������ǟ ٟh�z��!�3�E�W� i���������ïկ� v���/�A�S�e��� �������ѿ�������+�=�O�a�s�^���$UI_PANE�DATA 1��������  	�}/�frh/cgtp�/doubdev�1.stm fn�ame=FOC_prim�������"�)��G� � � fr/SpeedHelp��s߅��ߩ߻���)������ ���:�L�3�p�W�� �������� ���$�� ���  }m���|����v2��g.sh{t ��dual.��������w���Z� l�/ASe�� p�����  =$asZ�~���@� '��&��}�//*/ </N/`/��/ ���/ �/�/�/�/?r//?? S?e?L?�?p?�?�?�? �?�?O�?+O=O$OaO� ���E�à/�O�O �O�O�O�ORO#_�/G_ Y_k_}_�_�__�_�_ �_�_�_o1ooUo<o yo`o�o�o�o�o�o�o 	|O�O?Qcu� ��o�0_���� )�;�M��q�X���|� ��ˏ���֏�%�� I�0�m��f���( ٟ����!�3���W� i��������ïկ� N���/�A�(�e�L� �������������ܿ � �=ϰ����ϗ� �ϻ�����2��v�'� 9�K�]�o߁��ϥ߷� �����������5�� Y�@�}��v����� ��\�n��1�C�U�g� y������������� 	-��Q8u\ ������� )M_F����������/!/)�F/��5/r/�/�/ �/�/�/3/�/�/?�/ ?J?1?n?U?�?�?�? �?�?�?�?�?"O������$UI_PO�STYPE  ��� 	� .O�OTBQUI�CKMEN  �cKrO�OV@RESTORE 1���  �O���OS�O��m*_S_e_w_�_�_ >_�_�_�_�_o�_+o =oOoaoso_�o�o�o o�o�o'�oK ]o���H�� ����o�0�B�� }�������ŏh���� ��1�ԏU�g�y��� ��H�R���Ο@��� -�?�Q�c�������� ��ϯr����)�;� �H�Z�l�ޯ����˿ ݿￒ��%�7�I�[� m�ϑϣϵ����ϓGoSCRE�@?�Mu1sc�@Wu2�3�4�U5�6�7�8�TBUSER�����Sks�u�3u�4u�U5u�6u�7u�8u��T@NDO_CFG� �cK��T@P�DATE _��None�B�V�_INFO 1e��	�A0%�� $���S�6�w��l� �������������=�O�2�s��L��OFFSET ��M��t��@�������� ��'0]Tf�� j������#@,>��O�
y����UFRAME�  t�����R�TOL_ABRT8����ENB��?GRP 1��I�ACz  A�I# G!��G/Y/k/}/�/�/�/�+��@U(��+?MSK  %	����N�%�%�	PRT50_R�02��JVCCMf�����l2MR/"2�cI ���~��	��^�~XC�56 *�?�6g�����$�5~���A�@� p� �[> 	�H)Ot�JO\O��O�1�O�O"E�%A��|��O�O|� B���	Q|�U �O._uOR_!_v_a_�_ �_�_�_�_�_K_�_*o�o'o`o_�o�oi4I�SIONTMOU4�4����es3��σ�υ�0>! FR:�\�c\��A\�o �� MC�f�LOG�o   7UD1�fEX|��' B@ ��br3qZ�3q���t� �  �=	 1- n6  -��tƌ_rt�,�vDA�p=�����qt�2r>xTRAINI�r(�q|��s
~�d�i�3��; (Ma�uz� Amz���������Џ� ���*�<�N�`�r�Z�h_FpREv0�6)��2i4LEXEs3�̘;��1-��_>MPHASE  �����Pj3RTD_�FILTER 2]��; Ԋ�O e�w���������ѯ� ����
S�8�J�\�n����������ȿڿg6SoHIFT�"1��;/
 <o|%o5��b���9�r�I�[� ��ϑ��ϵ�����&߀���\�3�Eߒ�i��	LIVE/SN�AP]�vsflsiv������c� ��U����menu����|�A�S�*��s2�6*	@�?��hhcB@ �@@�9�A(�B8s`s`�CA������0�@͖�� ��4�7�MOs3���� ��$WAITDINGEND�h�([�O0��/y��j��S��v�T�IM5����G `�������������<��t�RELE�/�X��o #2Y�_AC�T�Т@2u�_�a ��8;  L_L�ATCH����R�DIS��/�$X�St2�6+�:�:B�_$ZABC/#���� ,H�PeO?�Z+IPs���Oo/� /2/�MPCF_�G 1�g 0�pb�z/@/MP��g1(��Mo�/pa8���/?�/3?�$?�7;M?7?!?�?�E?g?�?{?�?�?	a� �0OO!O7OEOoK��S �`�g��YL�IND5��g ��phd ,(  *�O�Mhc�O
_�O._] �?d_v_�^�O �__�_�_�_oH_)o ;oMo�_qoo�_�o�o��o�o o��#29�g� �p/^ n|�?����9N���7��A��DS�PHERE 2��M�eoA��o:�w�^� ���o�я�_o��� ��=�$�a�H������� ���ߟR�����9�`��]�o����ZZ� ǭ