��   #L�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG ��D�HCP_CTRL~.  0 7 �ABLE? $I�PUS�RETR�AT�$SET�HOST�  ��DNSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!MD�* �D $PRIM�AR_IG !$?ALTERN1��<WAIT_TI�A � |�FTޒ @� LOsG_8	�CMO>�$DNLD_F�I:�SUBDI�RCAP�  �q��8 . 4� �H�ADDRT�YP�H NGT1H����z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV�  D�P�INFO.  o $$$X�<�RCM+8 ?$| ��QSIZ�X�� �TATUSWMA�ILSERV �$PLAN� <�$LIN<$C�LU���<$TO��P$CC�&FR\�&�JEC�!�%�ENB � ALkAR�!B�TP��/3�V8 S��$�VAR79M ONx,6��,6APPL,6�PA� -5B +7PO�R��#_12AL�ERT�&�2URL� }�3ATT�AC��0ERR_oTHRO�3US�9�!�8R0CH- YD�MAXNS_�1;�1AMOD�2AAI� o 2A� (1A�PWD  � LA� �0�ND)ATR=YsFDELA�C2@<�'`AERSI�1Av�'RO�ICLK�HqMt0�'� XML+ �\3SGFRM�3T̑ XOU�3Z G_��COPc1V�3Q�'C�2-5R_AU��� � XRN1oUP=DXPCOU�!S�FO 3 
�$V~Wo�@YDU�MMY1�W2?��RDM*	� $�DISc d�S�MB�
"�BC�l@DCI2AI<&P6EXPS�!��PARQ#\�RCL^� <(C�0��SPTM
U� P�WR�h'g�Ro� l5��!�"%,�7YCC�% 0��fR�0�eP� _D�LV�(f��SN�IFF� � ��$?�s_ST6�$: GG�$0qd'v�PP�$�@^MvBUFF�&RP8bq��3IFI��>�XPOSAV�dNDп!\3� ��0WEsRUE%�EOWN���AEa0�d(ez$(�`o3 �o�b�X_`�#Z_INSDE,C%�OdpE�dkUR4�D����t��   t 9�!�`MON�m��D�n�HOU�#E�yAt���������LOsCA� Y$N�0oH_HE��P�I"/ 3 $A�RP�&�1vq�W9_~ wDEF'�;�FA�D�01#�HO�_� �R܂EL	%# P K  !�0�WOa` -pACCE� LV�k�2�q�K ICE��p ��H�$*�  ��������
��
䨐�`S$Q���  �:�$X'0 ј
���F�����ܐ���$.� 2�T!�����>���� ���!`������^���@��ί��������À_  �� �4�F�X�j�|��������Ŀֿ������ _�FL)p Й�� U�����������nx�2����SH^)`D 1�d Pᯤ�����Ͽ� �Ϸ����<���H�#� qߖ�Yߺ�}��ߡ�� ��&�����\���C� ��g���������"� ��F�	�j�-�c����� ������������ Af)�M�q� ����,�P t7�[m��� �/�:/�3/p/_/�/W/�/��PPP_�L�A1�x!�1.�"0�/{&�%1|?{&255.;5L�/}#���#2�/�
>o0?0?B?T?f63 p?
>�0�?�?�?�?f64�?
>_@O O2ODOf65`O
>�@�O�O�O�Of66�O
>OP�O_�"_4_�RC�G ��$���,��C�?� Q� �/�^<�_o1ooUogoyoLo�o�ox(P�o�o�o �o'9K]����^vw)�1��1��
ZDT ?Statuse��@�R�d�y'}iR�Connect:� irc��//alert�����ӏ �x�.��%�7�I�[��m�!��P�bb�d��r�����̟ޟ� ��&�8�J�\�n�����$$c962b�37a-1ac0�-eb2a-f1�c7-8c6eb�53b57e6  (�ӯ&���	���-�{%<Qb��X��R^��zP��Pc�
�Q��T,$�b��! ��ֿ������0�� T�;�xϊ�qϮϕ��π�������,�߀ ��Q�%�PDM_�Q�	�+�RSMB 
�)�Qd3&߀_������&��_CLNT �2�� 4�t ��"��|�U�4�F�� j�|�����������-��Q�c�B�����M�TP_CTRL ��%�����tQ� ��	}���1U�|���NIFF ��ߺPNONE�b�  fr�:sniff.c�ap�frs:�diss��.dg��Ë��t �v���Pm�Gaz��y����ԁ�z�6USTOM �m�|�$�P ��$�TTCPIP�g�m��x�U� TKEL�$�%�Q�{�H!T�$/�rj3_tpde� � R!KC�L,/�R}��E�!CRT�/y/�/�R�Z$!CONS��/�
@!smon�/Z$