��  	2g�A��*SYST�EM*��V8.3�382 5/9�/2018 A��  �����AAVM_WRK�_T  � �$EXPOSU�RE  $C�AMCLBDAT�@ $PS_ToRGVT��$X� aHZgD�ISfWgPgR�gLENS_CE/NT_X�Ygy�ORf   $CMP_GC_��UTNUMAPR�E_MAST_C�� 	�GRV�_M{$NEW���	STAT_�RUNARES_{ER�VTCP6J� aTC32:dXSM�&&��#END!ORGBK!SM��3�!UPD��AB�S; � P/  � $PARA��    d��ALRM_REwCOV�  � wALM"ENB���&ON&! MD�G/ 0 $?DEBUG1AI"�dR$3AO� TY�PE �9!_IF�� P $E�NABL@$L�� P d�#U�%Kvx!MA�$LI"��
� OG�f �d8�APPIN�FOEQ/  9�L A �!�%N�! H� �&�)�EQUIP 3�� NAMr ��'2_OVR�$�VERSI3 ��X� COUPLE�D� $!PP=_� CES0s!_81s! �L1> �!� � $S�OFT�T_ID�k2TOTAL_E�Qs $�0�0NO��2U SPI_IN�DE]�5Xk2SC_REEN_(4_27SIGE0_?q;��0PK_FI� 	$THKYGoPANE�4 � �DUMMY1d�DDd!OE4LA��AR�!R�	 � $TIT�!$I��N �Dd�DPd �Dc@�D5�F6�FU7�F8�F9�G0�G��GJA�E�GbA�E�G1B�G1�G �F�G2�B�)��ASBN_�CF>"
 8F CNV_J� ; �"�!�_CMNT�$�FLAGS]�C�HEC�8 � EL�LSETUP �� $HO30I�O�0� %�SMA�CRO�RREPR�X� D+�0��R{��T��AUTOB�ACKU�};DEVIC�CTI*0�� �0�#��`B�S$INT�ERVALO#IS�P_UNI�O`_�DO>f7uiFR_F�0AIN�1��x�1c�C_WAkd�a�jOFF_O0N.�DEL�hL� ?a8A�a1b?9a�`�C?��P�1E���bEX_CN}!� � �'$� _y �0Ya^aXsgOPTC1}bXI��PEE�xs� TOds�RE�cuvnx��R�yp_RDY_�OU�}IAL-uG�W. l @8 [p�0tt[p&U� �1�3B�� ��"; �o 0� uR�"SwCANM� �-u{POqA DF AVAILua�|�@�p��r�������-u, \�p�A>!RDINGByq.�COMR0T�pA��3S�PIR��A�E ADYs"MO<� �cE D [�M�c��B�REV��B�W� K0XI�� 5�R  �� OD�Pz��$NO^PM�;� p���/"��� L���� Hp��0D`S� p E R�D_yp{ ( FS�SBn&$CHKBoD_SE^eAG�q��"$SLOT_���2!�� V�d�%�哝3 ��a_E�D{p� � ��"��PS�`(4%�$EP�1�1$O�P�0�2�a��_O�K�UST1P_C�� ��dx�U �PLA�CI4!�Q͢��qb��M� ,0$D�ɦ��0�`h�EOWB o��BC`S�r�ra�(ra��_M�O�0����`���"Fp~�����PSWN#ȅ�3Z`EN 1SV�A.�K�D� Z�3UL� A� [�q�� ǱM! �R_LIMka�DI�`PU�P�"س߳�r�2���TRQ �S_BN-ORQ]6�U4a��G�_RM.őtP��3j�؀���5�CT1LĴ��%�LMñ/�b��I\�]��ST'� \���a�Ň�Y#�������BIGA�LLOW� (�K�"(2�0VAR�Մ@� ��BL8�0�p� ,Kva ��P4�� y p�X՗��CFٔ Xf� GRP0+�MB�`�NFLI��Ӈ0U��P&e$� SWIT�CHHvN�P؂r�_��G� �� WARNM�`#!W�qP�V�NST� ��-�0bFLTR��T�[��PT��� $A�CC1a1���7�rb��I�o"��RT�P�_SFgh@CHG*�0I���T-��1��I_�T� �r��K�� x?ppj"�Q��HDRBAJ; C�����3��U4��5��6��7��d ��9{2XPCO1� <F �ߔߦ؈#�92:�LLEC]�
"M��I�b�" ��1؎!9��0T_}R   4F <�Ft�=b�)2��oܴ�`T! |� Bx������P�_��TTiO���E)	EX�q�.�b��焺� 2� � ���"[0`Ay}Rf�����4���/� #D"/�g�Q06����L���A$��Bx�1P���M.�ܽP�# ��TR;IG��% d��8�P���`A����e�p�5���  �:�^�R��& t�F{LEE2$ANG AgpTBAO���1� ��!�Ӑ���0+�P[`%����'����m 2b��X!;���"J;�_R,�erC�r,J>�w(�,J�D !�Ҳ)�ݱ���0}"o�CP_�POF7�( @jP�ph�p���IT�c�pNOM�Px%3�S��B P`T) w@&�L�� ��PA���b RA]q�Î4�X��
$TF^�:D30�sSU�P�!���(c1H�u/`1�:ESq����û�WA�֜cAb3YNT��� DoBGDE7q*V;�P�tq��J�;�P�#AX����eT~��ÛUF� d3C
+� � EGY�PIV;�*c0P�GM�H�M�I8@�FF�GSI�MQSTO�a$wKEESPAT�Р���2���2����!L�64FIX
, ��v�!dC_� ��`RY�kSCI��hVPsCH�PhRADDdV��QqU�Q}W�Q�X;�_Pl"P_�P�f�Q� =��Rв�51]�3B��*CWE��-�p`XF� nVGc}UGc�V�Xpc�Me�Ypcgg��!MC��.��@�SM_JB�b��a�S�g� ��e X�b�/� �e�CHNS_wEMP��$G�0�w[��0;3�1_F�P;4�1TC1v~wT�1{��Ft�u �_V`
���lqi"uvJRS�~��SEGFRA=�ܱp�RSTy�LI�N���sPVF(���!�19D0��y��rl"�%��r bH�!G'1` +�/��#��q p(��q�`����9�jH��aSIZ�od��C�TN��0h����qR�F�!,�ms߱s{���p��Rp�pL~��0p�CRC����;�ఀ�p�1q��1r)�MINI�1qr!/�߁�D�Զ�c�Cr��� �et���w����EVD����FÑ9�fsFVp�N� �a�ց��;��<c1�30�1V�SCA��0AQ��r�r1^�
2 ����t?��RGР�"?�Fțpl�FqDߵEqLEWZĮ S�����/��p�
�v�3� �I�[���P�E��R�	0HANC~�$L�G���A$YPNYD���ARcPN��`�q����Yse�ME%Q0�f��@`�RA��e�CAZ$p�����5Oz�GFCT��Π��F��pL�Fp�`� ADI�OȆ��������0�������SGw#���BMP�t���Tq1AES�Pœ���|��H44  	��I���CSF5��$��YC���`���d6� ;5$��SUP���ARM֢ւ��=pS@`.A �<Q�KP�#�#֝�#�O+�O9�F*+�F9�N+�N9��'���V_���DKI��DK4s��SUL�9���,�DD�3��GUA:�R��R��R��T�,�R��R��S�0\���OOR��U�p � -�q��|�{�|���|�Q|殣UTOOLw���������� ����⮣%�-؅�%���%�U �M`"՟�]ҩXWu]�YO�ZO�NUk�Vk�WO�I�����X�`H!
7 x�؀��$AT���7�CZ�Nqp�qI�MG_HEIGH��A��WID%P�qV�T$pAC���9AAp_p(���T�EXP#��D� �CUPMM�ENU�8�TI�T1$PRO�G_UD%W!�q0BZ�_~���9��UU ��Ax�6NO��ADE�����ޯ3�p7���APn�d:����� d��AERR9LV A ; \�0���OR d0_IDx `�0�pUN_O\�>��$SYST�UIǱS EV�3�paTPXW)O��A <��Ke1�B� �T �TR�L@= �U AC��p�4��INDˀD=J\TLAY_R��A��"��PL a�bWA���ESE�RVED�'!a����"�UMMY9�R4"10RC0DBd��@>�«APR�� 
�DPOsS_~@@? F`�-Ӆ���Ll)@Ly/#�X�8�A A�/^#���PC@B�/~#�H�PENE�0�Ts�C�/�#M RsECi�@DH��Cm  ?$L/3@$l#�B��@;�p�W��rN_D1��@R	O�P�qT�?�r�8� >@RIGk�6�PAUS�3�tET�URN�2N�MR_��0TUx0�^0E�WM�r�QGNAL<}p�B$LASˁ�3�&qA$P�B3$PѰ9�C@�cPCD��8�DO�p��Y4E12�_6GO_oAWAYo2MO�q�!�g���DCS�S_CNSTCY4`E L(�0;p[妉BID-ѕB2�J2
�FN7@O\�2iuB�ѐIj0 F P7 $Z�RBV��S�PI�GPO XI_#BYɢSWT��tC�HNDG�!G �H� ��Gap$DSBLIO�VeT�F�^Y� tCLS�aH�FR8 OUTzYFB�\��FEi1Z��S�D4tC��IFRDOq%�^�MCpd�P]b��R��H�W ��D ���uBELE��J �T�@�0سINK_�N��`bZ����FHAX�Fj�ր$q A悏  �tC�A�`K� ��MDLIb ?2J 
$�p�P��#��c2uC�k�c2u�cJ�cւt2r �} )tw�PdrE	�BZ�{�tCSLAVs�L�rINP�PV�P�~ytA��M� %$���= سV fV ,֥FIM�ro��sID2�s��vW����rNTV糺rV9E��tSKI׳D�H���9�2i��J��x�� ��SAFE�f�w�_SV�EXC�LU�E��ON	L� ��Y�TD���.bI_V0���PPkLY R��HIr���v˃_M8��@VORFY_�ɂMȣB��O�����1��d+�U�O�@΅LS�0�mR=$36RP��SW$SE�P{$zDb!�P��q�A`�s����Q N0��T�A�� C ���D�u�O�B�@Y��tkVL�FR�B������B��TCd\�"P� D $ �BA�Y`_cB�!�IpK�_��V���V� �X�rv��K�@QE�'RG:�0��`�P   H�rS}GҠ R ��`CUR�0�1��ʢq ���1@wϨvߦ��UN� mT��Eʠ8dE�0K�'�$�;�,�H�O � I�"�S @� F	�K	$TOT�0�C=$ѤZ�:'4F"d�MPN�I�"T�B�����A�-�ԴDAY4LOCAD�D2$��3#5Ro��EF��XI�R%U0(!�O��a����_RTRQ�5�V:�� =>�ErBJ�E��T���`U�`�"�:��DX�A8� .�5�W 0A�����c9p��;CM0oSU��0����CAMp 3Xr�� NS����IDL��W���S�V�GV_���`����DIAG��5�Y�p .$V�0SE(�TACJ�Hq>� E�D� GrR�"�EtV� �SW{ѷ1K����29��`�VIp9�OHOū�PLݐEtIRfGrB� �¨Ï�2FqB���B�����p�����F���`X�`>�z@B�RQDW&��MSB�>�A� ��<i�EtLIFE�J�Y�D!TrN{�E҄�$�$y�E�C�W#�Cn@H��d@N�0Y� �1FLA��#�OVn0�� |�0GrSUPPO�lQTr�_��ե��C_X�^A�Z��W�nA���$XgZ_Ab"HqY2i�ECn Tvw0C�N� �AԈ�CT�tZ� `�@CACHE�Ͷ��cץ���2SoUFFI��p���2$�3#b� �L�DMSW��[� 8<�KEYIMAG�3TMC1�1ૢ-|r�1AbN_D���A5�\� $[CM� �[�BD�Q<!\MAC�2�PD�1�\�A��Ĕ�P_OF0T2��Q�	ST��� �MSG�
��b ��1�nArP\2� M�1�VN� ��DV��PRDC@Nz�����\|pFx1>�ANLGF�[P�1��P�A�A�ȕ�b���7c�fpOC�VIE��$1] ��aBGL�$��s?��|�\�D��^�:�1`STE�! T"&@\$��\$��\$�\ EMAI�`�1ݱ�d�eQ_FAUL���_$"�3ݲQ�j@U�'�T�%LTT�  /` dƱI4�  R�y�&2�rP�&fc�'�(��'I�,Ђ �!T�REђa< �$>3eS����IT5�BUF���q���D9N���SUBj4�D�C�t��?2�DTSAV�5w2?Ј򼁏���7��(�P�4eOR	D��� _j0�5ΰIGOTT�����P�aM�u;D��8GAX��e��Xj0��3_G�{�
��DYN_D����b��� l�DU���M����� Iƹ���P8��c�� � ,��"CC_R��IK���Bࢄ�DopR)�E�(�AD�SPA�BP�`-YI�M�3"SHQ�c�C2�U��G����CM� IP���C��D� "STH����SR�T�"SH�SD%1"SABSC'�����V�d�V�P���T_DfcCONV���Gfc�T��Vj0F�{�TpdS� _A��SqC$Ҁe�CMERĄ>�AFBCMPă�@�ET����dFU��DU^0$���E�P҂CDY�P,@�#� � NOAUTO��e:��dε�d��PS�eC��e��Tp�  ��d?@��f/H *�aL�p�#%sLgF�{�E�Ct�� Av��Av��Av�Avb�(Av!Av8>y9>z{�T@xJz1Wz1dz1qzU1~z1�z1�z1�z�1�z2�z2J{Wz2�dz�Nw~z"Nw�z2��z2�z3�z3Jz3W{dz3qz3~za�[w��z3�z3�z4�r �t���UTP 5�g� � $��MeI�NLfPLCWAR�MS%�� >tRL���FKAC��S����Pj�1̚2���q�r���Jq 5d�EX:E�Bh <H��(�� ��� Me�@6��e��FDR$�7iTJ0VE��4Ap~�t��R~�REMM�9FVq��OVM�C���A��TROV��DT�0êMXҬ��_�8��ª!�IND᠎��
�%0~�$DG@jA��̠J ��j�DNƎ̠RIV|`���G�EAR�AIOa�K����N� ���_�`x���Z_MCMn~�L�F��UR|b�j ,�a�1?� ��]P?߰z�?߱E���W�1�Y`i�k )�PRA61�RI�% ��5�7UP2� l qpv3TD�P52?į ��M��G�  �+�BAC�Bm TR w2�0/p)$PROG���%�`�Bq���IF�I����Y`*pw��Px��TpFMR2f�n s��`qBt�L���x������P��Q��哢_�qK��LIMI� ���dC�_LvW�i�<�CL�F��DGDY��L�D��;�5��2�������G%o� J�� T�FS@H$p� P%�&���+ ~��$EXI� >�&�1P^@`��'�3_�5_�s�G�Q��q ���ybSW�5ON��D�EBUGJs�☥GuR�U@cBKUK`�O1� ~�P�O.�����k`����M�SZ�OORC�SMzZ�E�2  �������_E r �/P70IM �TE�RM/�s8�ZB�O�ORI��3�t8�.� �SMyOw24�=u8�[��c w��v��UP"w�s -����r$D�ʽ�sȐG����EL�TO�!$USE�pNFIG����ʰ�� ]���t$UFR��$�`��! ̗ee�OT.`TA��P��@NSTa�P�AT�QTPTH	J�Q�`EJ �2����ART�0�����1�"���REL�
yASH�F���\�_SH�ORx`�cu� ��$��� v��u�OVR�]SyBSHI� ��Uz�b ��AYLOwPrA�AIXa�\�P�f�PERVIp'�P�
 �<a�Jq������RC��eASY1M�A�e��WJ�����EÆ�c�aU��a��A��!�e�P�[SDaORa�MF��̆����x�"�����  qA\�sHO�+�y �B�����TOC��|�ᰱ$OP� D`,P/sya�0��O,ա�0RE� RcyAXp��3]e� RZ��%�(���e$PW�RP�IM�%XR_�#VISv�o��UD�s" �z;�$H��!^i0ADDR6�H!�AG^�1w1p1k�Rj@\0@�{ H%�SF` �1Js�5�5ds�5qsxɑ�1l��HS�`�MN�| �`�`�"�Q�SOL�xS�@��E��f�AC�RO0��!ND_�CxS�bV54aROSUP@ch"_
PIxP�!i!1=�҅CK��I Jp�I���Hdp�Iqp�Il~p�AC�IOAc�AVED�G�C�ED<�3��} $�� �_D������2PR�M_~B t�_HTTP_�`H��~ (�`OBJE�^ar04$6�LErMOS� �}��2H�a_�T�RS|Ր�SDBGLV�R�$KRL9HIT�COU����G�pL�O�1�STEMP��S�RԢ� ��� SS��NdJQUERY�_FLAEB�HW��q�����0 I�NCPUB?0IO Rf�QItib�4ja�4ja�qr��IA_CH�KCM�P �8#p+q���PxV�RМ��pNTL�2�aR_t!~@�a�f A��7��R�h��_J��
sSl�QvIDzVA� p@03��9��Es-vEs<u�`PRp�a�r B�1�b�q3�yTrH�Ӑ�t-uSRP�~���t�wOPw�t����c�����W�`��ĒOT�Hm�N�$WA�z�!�AF�1e$�BF����aWT_P��cr�9RIv�I]��TYAZ Dp�qaU}R��R_BICL�BYPASv�A�b@m����R�`��v��Ӱ�$Lh$�
$F����C
  \|߃�P � 8%���X��{rMATGRIX�bC�*L� :3 �aFEL���0G� dE�-�O�K/��~P�6�SHA��I�ZP�ATA��$7LNT�CH#e����^C )�d�cP�1� 0հh� 2��V"l@
PD��!9հ�(  dc��1� �-��h�� D��v�����:���ROB �F��^P镇��U@��8�SL����CAkLI�b�&�DO?��o��4�a3P;OS�1�  =�-�BA��ف! cP��b����1�T X�$BIA!3�a T��@�aK�����2�2�9җ�j���# _HAN	� Q�Рj����S�@#2�=���j��*;A�X$aOA�yU�RAN��Ax{rH�X@S�b��_B;P�B�!�q�����UBP�R��q��O��"��E�LBOW�a
� �
̕aL+��G� ���ɱM��x�p�3Y�SLICM0�)��#5E�r��P8XP#0��OSG2Ph�YSWAR$�"H��t!��h���W��CH Nx� w�)�ESsYN��zSR_fAfJ�H_�pI�ES]a�
X�R��IDLL�a�cUN��S&�`�݄����WNO��D��'@O���a��R��)R
p�_��LR��5@��'����P�2 q 8o�R�w��Y��o�L@�~@v�{��බ�@ARGI��L_	N2P �A���a�g�o�d|�R���බ�1�� .���V⻅��鲟��LA@�sM��a��� tؑ���w���  ��P��OT&���22F �������*!PgQ��2�MtW���t��PAI��� � x�@t"RBâ�!��	}d�Yt'|�EY�s_|���B	J��v������t5 ��REAI���便1v��咾HE7R %a�� ����֓Π����}򝴓 ���^@UN!�� S�RM؃>�XpJ�J�(�ECKC <��`��0�Sr�A�r���_T�a ����2���0ݑ��2��0R#EF5�q�2��10,�3��0ゔ��D<�!�qETHO��;1����`Õ�W���$�B�Wh@(�IOL�\0C���ܑ�WT������r�f�$C���"W��f��WTP����� '�c̃TF`B��ʃ'�WaMYD {r���s�$B6�P)C c�xu���c���l7Vp��1]~�y���$FR�`0{�`0W' ��1 5�v4�u7��~�@4��?;vW�pI}62��2�6��2uuW��"�WT2_	�FH&A� TyƯw;$����v�� 	<����	�Rt^��j�����IC3[D_s��(��oTPGLU�AD����BINI�VOX�!�D�@AZ͡��W���8pߤΣ3�z��1ׅz�2*W1_P�1�G@Q2E[3EX2�B[nPSYnPbY'QPTn`�U��W�@�S@nP�W�Q�V�Q�V1T��2S�VEXTRA�1��b2���D$�G� ���N�@JR�\�3�PPEe@De �T-�FL㳽��Z�����y`PAųtdMEM^�tdP�oiG��C��a���BZT�@�P�a-��U��
�3���AP�� ��O���@[d�I��@� ����A{a�� �x�C0^`CN���N�C�SIV/�:�S� ���qH&�qJ��g�Q�`�p��
�j Qr�`�'� �aECf����f��U3�6@VERAT���#*�����	�D�LENF�H���V�ZS�MGQ�|�a�|�p�R��X2���Y��Z:rTOT��B���`� �B��a����{
�8:�uL�� 4�� �g����!�E+p� �CDPf�t �$`���MjhERG�q��Vd<�C�|c0���Gķ�Z䩕��E ϒ�!�ߑ�!�!�bQ�GS��}��a��p��INO�9�&�>�^p�N_XY�Id
g�Zn�Gv���&��� 2�C����Pb��]��e�l@)�P�$ANALY5w�b'��Q��_�Uu��b�I�c�� :a�Df�'�1��p� �  ���G��z�Up�R3z�А������I�^�BGD�� � �d �P��FIO�V�-�c'�&�>�܊�TAImsBUFEX�� �߲�ǧ |*`�}�MEֽ�a�Ir�SV�q�SV~�COq�On~�PATJ�)ex�dk� ��Be@�BOX�� @ Ҭ���_����ʁ�����^ ��^ �  �dݱ_��� �@�M|��p0�$ACTC�N��UPDi�A�l.Ҏ�D� �!0Н�D�Z�*�:tOM��$TE� ��aeq�ҭ��FL��a�N �a�v� A��h�3�  �u�"�v��\�>@�@��� VRWRT:�L�NTK*�ARCT�OOL�A`Ѹv�Z�'�_ � ` $ZPR1���B��TOK��џ���p0���'����R#VE�����.�W�1�@"���#PAP�ҧ
$F���D.�S�I�B���e�"��B�9 4�"�\߬�ALC�PEQ�j OLNK����`���Hq��K!� ��_��H@��Pq���u�_SLAVE{��b������������� �u�_�AS�A� T��Lq�&�fd$�p�RT� 	1�����~pH�5\P) r�U�{����n6^ >x^ G�TRTPK# ����G��
r磾3q � X��I�PAD���_NE�!��LAG�!� 5 ��#�q����d$FOCUS���Mq�TEM_AC�r�S l�� M�L0p$�p�NL7�F	 {GELA�!{E�F�4�$H8!�REP`��rI�ـ��b"Z�n��N��>��IRCA0"b�� � | v�I/NCYC�A8/!�M�3-@3CL'I��G<6�cDAY_��NTku��'��u�ΐ'SCAd �'CL'EAR�!�R��q@�P����r%5N_PERC�B �~!�@��C>C�7� r�p��1_OF�(>>�3�  G�qP� $w6Q2w�LABـ�2��7U��B7H�@xuHT ? ��UJR*Q{�� � F��D�~c0@`W�2˦J7*P�c�$J8I7_AHI�E4G7�6@8KI�AAPHI�`Q�#ChGDSB_J7�J8��BL_KE�a����KARE�LM� ��XmR ON�WA���_VAV��r��1EDAp�ty,НBq�rrc�Vs��@CTR����B	,�LD{�Ǽ x`p	��uNTaD�!TdT�L�ORQc^M�NTMO\VT%��PD��S2 RO�J�VTOms����;LG.T� ��э�B�W��p�`V�WcMR�W �VFD�XAI�X�X���V�XP]�U�PMOD�VRf�P�Rf Rf`RfC`RgX#_Rӱ���p~��O��LNA�2����DE����иa"pU��a�L�c�bwDAU�eEAD�a�I�r�`GH�s ��� BOOz�g� C/� IT�s�5tT +RE�pLxS'CRN��+Dr��� @�RGI����|@��#U��u5�S�1�"W�t�d#JG=M�wMNCH����FN�B�vK	�PR�G�UF�D��F�WD�HLL�STP�V���<p�;RS��HELh�D� C�4b�Ec��0�w��UF&��w���w�P8�G�y�PO �g�wub�Mɇ:��EXTUI�I 7`&3+ 7a�r���s��`���Ѱ���	��iuѱipNwQP����TAV=��T�%PUD�CS� ������O�!�O-�Sf#K�8�SD��xIGN�P����p��ѯs�DEV���LLRQ/��|���@�T͒H��U�8$VISI�T�b�A ��@-�oP��P��;�1�2��3'�EP��� � �)��T��Ku����1&LO�Lt4A�STo Rp��Ѱ>�� �$�в�C��@FF��Ҷ�P��� L��>R` S����Y�2��8��hs_ ��s0$��������{MC�b� � �CLDPo PUTRQLI�1RS�0�ɃăFL@���1���!D�A��R��D�šķ�ORG�0�����������3�фt��3ƃ �8P�Ļ��ķ�SOV_PT����	���p�x�RCLMCІ��(ߘ�4v� ��MFRQq�� � !)HRS_RU����!@ 0��k��`>�$���WOVER�c
M���6P�EFI��%�W ���C�� 1\�0
�4D$M�j1f4?8P�!PS� �	�sP��i����U0ABP?( }	�0�MISC�5'� d�aS�Rn��2LPB�p� ��q��AXPR�@��EoXCES8 �@R��M� {��'P��PT@��SC� O� H=1��_n0@��S ���/�L�Kra�y�;T��v"B_�@�FLIC�BVpQ�UIREɃvP��O|���VOB�ML-�Mq� [�Dq6 �$R:S��ڬ�MN.R��1��b�bX�uDCb��dINAUTyq�d�P@�p��N`RRa߃[!pbPwSTL�1� 4=07LOCV�RI&0V�;EX�ANGV���� �R`A���b���2�0��MFR e<�|�,�6�b�`���SUP2� \w�FX��IGGHq � �8P,�Ra �$-�ӆ,��@[⡲� ��������=�k1ܧ�@1�"P N ڠI�N��� t*MD'!�2)5&\�@$��='1HA@$DI�!@$ANSW�q@$ �p�Z@%D	s) s�O�3�n��0� ^�CU��PV~ �����&6 LOp�0�\��$&��P�&�2ո"�&��#�w��MRR}2�5�� �!��aAu� d$C'ALI��SeG�,7�2�RIN�/4<;$R:0SW0��j3�*�ABC;D_J�2SE���4!_Ju3�6
�21SP�@$=���P�4�=3�=�!CP���5J*��57Қm�O��IM*���CSKP��$D�`DS$D	J����Q$LUE;EUEKG _AZt��1�A�EL���2��OCMaPyт��`RT�a��C�%1��@�%v�1���H���JZ�DSM�G�� ���INT	E����׸"U�r���8Q��_�� �0$U?R���� P;Uw���IYDI�A[Q���DH?�>Pk��c$V90�v�$���$�@ ���$�Y�X1���H? �$BEL�@��}C.�ACCEL\���X*��PIRC_5R��`NT�ဳ�$PS?���L  �P)f��Pg�a�fPATH�Ybgc"bg31b�B�_��R��`�a���Q_MG���DD�a`xr$FWs� �S�ec�R��hDE�kPPAB�N9gROTSPE�E�b� S�KA�D�EF���Q1`$U�SE_80��P$�CD���Yp�Ps� ��YN��A<@�v@W!n�qMOU�aNG��`OLRc�tINC �$�b�d��wA�ENCS80���)aX�R�&`IN��I1b0� ��K@VE�p032�23_U&A�D�/LOWLP��� S��ud�D������P�1��u��C/P+�MOS}���MO���s�PERCH  �� 0�h�̀ĆV�΃�g� ����G�Bjup`d�C	A1b#�LڔC��G�,��g�b�}�TRKׄN�AY�#��� 1b����	�F���r��MOM�r��н ���c,7��dc�0�DU@�bS_BC?KLSH_C1b$� �p��1��s��C��rM�<�qMECLAL۠*�p\�Ӑ��CHKS�:e�S�pRTY��!"�ޥ��!_����'_UM��ϩCܣ�a�SCL���LMT�0_LРC�g!�E�)���e$�h��08��q.�j��PC�ԁ�H3� �eҥC̔�7�XT�P�gCN�_G2N��ɶ*�SF�Q��Vjr"���Q���1bŢ�CATٮSH��G2�d�v����`�%2a�)�@�`PA٤&�r_Pإ��_(@�������Sѩ��Ĭ�JG0e�U��R�OG�� �TORQU\p�5������`����` �_W땒��A�Q?ԨS>ՠ�S>�Y�e�T�I�SF���1��2��A�`VC"�P0�����1��Q�8�����JRK������ֱ DBL_SMt�q=�M� _DL�Q=�GRVE�>�S>��S�H_�#�e`l��COSy�@y�LN ���գ�P���@�� p�������Z�୆��MY�����TH|��9�THET0m�NK23�Sc�S��[CBh�CB�SC��S !��pԛ�S��h��SB�S��s�GTS-A8qC�1�G���G<����$DU��F��,2�q��$AV�Q��$NE*DsI��ຣ�ITW$�PW�A�[���k�v�v�LP!Hy�b<�bS��� �����b����
���PV�V��P�V��
V�V�V�V*VV H�����B���H�H��HHH OJ�O�OQ)�O�
UO�O�O�OOO�Fb���)����$�SPBAL�ANCE�4��LE6��H_[�SPQ���<2��<2��PFUL�C@8g2O7g2��)Z1=��AUTO_�����T1T2�9�R2N ���R4��4WQ̑i0G (8b�S�TS�O�@�Q>/�INSEG�R���REV�6��%�DI�F|�NY1�3GzR1ل@OB)Ao�H����2
�4���'�LCHgWARr�RAB��~��$MECH��(�q�A��AX��P�M��F}�R P� 
p�B��Q�ROB���CR1bU�� ���C�Q_��T �� x $WEgIGH�pm�$�d:S��I�qb�IFTqN�`LAGrl�Sr�@rBILsUOD�Ր��QRST�PQRPAo�RP��P,�!Q*P��.P
�p�R�q�� � 2ܔ�VVDEB�UbSLZ`�R M'MY9!e@Nu�d�m�$DZaށ$��P��J� 8��DO_`A)Q� <=P�V�0���qN�IB�R�PN(�_h_k��p��RO|� �/� "�T����T*A�T$`TICYKcSw@T1,`%�c���`N���0Sc��R�:��q�B�e�B�e3`P�ROMP�sE<B $IR Ќq��8r6�UrMAI$��q4�r/u_mP-s6@t���pR3�COD�SsFU�p_VID_ր�qu@r0G_SU;FFp� gS�q6q�bDO�g@�e �P�g�y�u�B�uѯt�3d�P�=PH]@_F�I�Q9�ORD��Q 0P�R3�����q,`�Q6e��4 *FAL_NA�haIpW��eDEF_Ig�W��fs��e�R�f��T�f���e���fIS�K ��Ka�0�d��c�q���T4ұd��RDP�0���SD��O0>JbLOCKEu��s��o�o�g聯r�pUM �uW��t���t���t� �r���u���t���r�V ���s�@&Q�uW��u@���s�-��x�`P[@ ք�`�` $`Wh�g����W���QGR�K  � h �$���2TbX�`TM�Q���^��bf���]cE�R'@TG�F��� ��Q�*P� � o$GR� S�ID��B�6�#�\��Ip6�R�3�b ���sS��a/���.�_�9 ^@>�R�!���H�MSK_�0��� P=Q1_USER�1�ұ�pv@����1VELV� ��v@ٲ͵�AI?��0��MT�aC�Ш��  �`;@R�W��RE(Pg`��OPsWOਰ�, `�SYSBUtJ�S�OPA���I�TL�U�K�6@P����r�PA`���téBJ�OP�pU(�f�[A�R�Q��OIMAG&��0��f�IM����IN/������RGOVRDDb�Ű��P�����@��0�"�ծBL\�B�T�2�PMC_EQD%`�@�QNt MD�t�Q�R1�R1<����SLZ0���.P$�OVSL�6S\�D�EX�����? laFF_��VR���p������p���׻��RR�`h�@pTU��� G@ z����EOypRIap~
�Ep�*�� ��8AE9CY���� H=Q�@��PATUS�
aC,L ��DXb�B��o�X����QD�BШ�� DAa����b�}s`c���Ї��XEi� $����������>P�h�UPR���܁PX�p����T2���X��PG�� $SUBW��E��W��+�JMPWAIT���o�LOW�BF�aM`q�ARCVF�=q�`�Br�RE��F|A�aC_CTRO ��c��IGNR_P�L+�DBTB�PP����ABW]p�� �Ut`��IG���`�1�@�TNLN��RT~'�NOMOTN�`<�2 �ERVE��Gؠ�A�r�SP�0 � L=P�@r�g B�tUNOP2�s �R��2DLY<��0a��J��PH_PK�T���RETGRIE+�$§���"pFI�� �x0P� � 2���DBGLV��LO�GSIZ�A&��K%T��U#�,D�� 3_Tl0�BMMh0�� BEM;RLP��F�CHECK I�%s�P����� 0��aA,0I�NX0K�ElPJ��R��PIP����$AR�dr����I�OR~+�FORMAT�Q ��R�D	$��UX0���J`�PL|vp��  O��SWIx@E#d�M�AX��]pAL_ �� $qAV�B^7�$CCV�D����U��J3Du(�{ Tx�PDCK0�|߂J�CO_J3&pPH�#�#2W��/�-�pPi0 .� �� ���PAYLOYA�#$4_1+:2+3w J3AR��J875�[6F3��RTIA4�u95u96V�M�PN�T�3�3�3�3�3�`B��AD�3�6�3�6�3PUB�`R�4�5�3��5�2��M"���� L$PI�D*&3@aA05L.7��.7ZCJ�pnJ^KIlCR0'1��F%�F2�Q/���
�SPEED�G i"�D��d�Fd���� ���FS�H��Y���SAMP�QgaTX�G�YS��MOV_�R �Q�P��Ͳ�T�%�Vr�80�YF0ͲR [�z4�Us ٰ��U�p �[s <S�X
k�T���Z�0hd0kPkGAMM��USk��GET�I�FI�vp3�
�$z IBR
�(I$c ��R�_��q�$��fE� �hA�n�`�fLW�mv|�i1v��f2�F y!C��C�HK��=��.I_;P ��R$9(a��U�w�3�t�6�yw# ��$�( 1��pI)�RCH_�D��[�܀��|�LE@ٱ���&�8�p�+ _MSWFL��Mk07SCR�75��T3#�z��W蠁0�Y��|� ����$$C� =S�����΁Ő�Ő À�SI�!�͆ـ��:�� VMz�K �2 ΅� 0  �5�Ձ#�/� �R� R�	u�f���ŐBπ�w�������e� ؝�t���1�9���sBS蠌� 1�� <� ~�������Ưد��� � �2�D�V�h�z��� ����¿Կ���
�� .�@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖߨߺ��� ������&�8�J�\��n���I�Q`(`LMT逕��b�n ��CIN����� _�������v��@��Z��΁��Lp0!V �Ή��G�LMDG� 
����LM_IF 
� ���������������+=N, 
m�u��B������>�NGTOL � Z��A   �$��P�FO U� |�Wi{�ւ a�� ҂���
/�/@/@*/d/N/t/�/$��� �/�/�/�/? ?2?D?@V?h?z?�?�?A�P@7CAT�?΅����b Sp�otTool+ ��8 
V8.3�3P/05#�4R�IN
1041�22�2�5IO �
F0'AJ "�
90BI\t�p�?s�AD �7DDE�0�9����GM Gl�obal 4 R�ev0� A�FRA�?�1J|D�6O`TI�V���3���CUT/OMOD�Y���P_CHGAPOcNL�O݁QOU[P�D 1
�� �IPM___q_�:_CU�REQ 1
�  ��H{\g��_q�����Sӂق �^	�1 Wel���SW]�s��SW}`K'fHKY �_͘�_�_to�_Pobo��o�o�^c��Handling�dH�ULR�jHT;a1�o�o�o��o�oB}c��DispensMeuDI2E'dL/hL;oI[m��� 	�'�-�?�Q�c�u��� ����������#� )�;�M�_�q������� ���ݟ���%�7� I�[�m��������� ٯ����!�3�E�W� i�{��������տ� ����/�A�S�e�w� �ϛϭ��������� �+�=�O�a�s߅ߗ� �����������'� 9�K�]�o������ ��������#�5�G� Y�k�}����������U�TO� �O�CDO_CLEAN_
TP�NM   {_������^DSPDRYRW&�UHI�@z@�R dv��������//*/�XMAX��07�A�a�AC&X�7�qDR�q�BPLU�GG7P8DS@�#RUC	Bx |A�3/�"O�"$SEGFP2`�/51x �R?d?v?�?�?�/1LAP/B>�s�? O O$O6OHOZOlO~O�O�O�O�OSTOTA�Lj&@V�UUSE+NU/0<[ �e`�!_�b�PRGDIS�PMMC2`�QCL1Z!@@$<TO-�O&58S_STR�ING 1	[
_�MPS�J�
NotAtP�erch�VIs�ItSaf�t�R�CycleInt�erup�TPr�oduction�StatusFP�Chut�X�Q  n�Mo%o7oIo[omo o�o�o�o�o�o�o�o��XI/O SIGNAL�UHPFr?_ITEM1%# q������� ��%�7�I�[�m���������V3�[3 [y͏��+�=�O�a� s���������͟ߟ���'�9�K�]�߃WOR0�[����c��� ïկ�����/�A� S�e�w���������ѿ8����PO�[FP	-����P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ�(�DEV0���DϾ� ��
��.�@�R�d�v� ��������������*�<�N�PALT�u�O������� ������	-?Q cu������c�GRIM �[�� �ASew��� ����//+/=/@O/a/s/�/�@R� �!1�/�/�/	??-? ??Q?c?u?�?�?�?�?��?�?�?OO)O�/PREGy�b@�/;O�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_��_�_/}�$ARG�_��D ?	����a�  	$/vW	[$h]$g�/w�Ei`SBN_CONFIG 
k�;qWgCII_S�AVE  /t��ayb`TCELL�SETUP �j%HOME_�IO/}/|%MO�V_�a�o�oREP��,* _;q`UT�OBACK�`�mnFRA:\�OK ,OF�`'�`��OGzx� �~ FhOM���
���@�st���F�n���������ȏ OE[����*�<�N� ُr���������̟ޟ i���&�8�J�\�� ��������ȯگ��!ׁ  fq_Is_\�ATBCKCTL�.TMP DATE.Dx�4�F�X�j���ZFpEXcb �iaE�� A~�sCz  B�{�e|e��GRP 3�e�` 9l�{OC,<�OD�aOI�e8�J�йCܼ�����"�H����X�PORT ���	yra���A��OL�e�+�E��y���WRK ߻�ߎv��C��yc��.��INIx��uuf~CsMESSAG�`�#�a`wc5�ODE_D�`�fue��\��OVc���PAUS�POS !�k� (7�����(O�������� :�(�^�L�n�p���������U�P��TSK�  �ְ�z�FpR?CV_ENB�`mm���UPDT\�!�dys r�XWZDC8#�qj|STA �a�saXISc`UN�T 2I�c ��V���� ?`�������& ���h��J�"� 5�� -SS (��  �R $�#gS�3G�?��� ~�<�W�z ������]0�!~b�|d��*��W�ME�T� 2�PV�I�s�I��I���I���I��CI슠��?�M?�{E�?��?��>�^�?����SCRDCFGW 1߹�p��e�b�{/�/�/�/�/ �/sOJ&�c/ ?2?D? V?h?z?�/�?~�?�?��?�?OO*O�?�$IqGR� g ��`C�kNA�`k	Itn]F_ED�1l˿
 �%-�EDT-NOz�O__p/j �e-Is�O���_q���G�O~_ ����E2- hg �_p�L_q1�c[��%	PRT20�PICK�_�m
 ��Z�P�_
nP_�g�V�@o�_oP3?o{�Q12�_�l�]ho�o o,o�oPo�C4�k �of��"U4��o�o��C5�G$�k }~ �k���Z���C6�����7�}~̏7� ~���&����C7o�ߏ ���}~���J�\�򟄀��C8;��O���o ~}d�ϯ�(���L��C!9�w�T���~}0�����������ACR r_���1�����eϬ�о�T��`@CE!p������� ������!���mP_GR�P 3�� X�+�n�\ߒ߀߶� ������������4�"� ��P�$�r�H�Z��� ���������8�J� ��n�����(������� ������4"XF h�������� z0��:<f �Z������/ />/,/b/P/r/t/�/ �/�/�/FX�/�/�/ ?^?�/�?0?�?|?�? x?�?��?$O6OHO�? lOZO�O~O�O�O�O�O �O_�O2_�?X_,_z_ P_b_�__�_�_�_�_ o�_@oRoOvo�o�o 0o�o�o�o�o�o <*`Np��_o ������8�� �B�D�n���boȏڏ �����"��F�4�j� X�z�|���ğ���N� `������f�ԟ�� 8�����ү������� ,�>�P��t�b����� ��ο������:� ��`�4ς�X�jϸ�&� ���ϜϮ�$���H�Z� �~ߐߢ�8߲ߴ��� ���� ��D�2�h�V� x���������� ���@��� �J�L�v����j��������$�BCK_NO_D�EL   +��/ G�E_UNUSEN�D(:IGALL�OW 1��3�  (*S�YSTEM*L�	$SERV_G�RPLL{ POS7REG�$��
��NUM�
���PMU' �L�AYER� PMPALT�_CYC10
 �	AULSU`��� �LW~�BOXORI��CUR_}�PoMCNV�}�101�T4DLSIBt���4, L��3/E/W/i/{/�/�/�/�- LAL_?OUT j	7 �r�9WD_ABO�R"K 3ITR�_RTN w L��3	 0NONSTO� K4 38CE_�RIA_IH K5��07~0FCFoG < �/� �1_PARA�MGP 1;".��?O#O5O��9C�  TN��W C�j@�V@�j@U�j@�V@�j@�j@��  D@ D��@	� D� D�@ND}A�MU�@�@�@�@U�@'�@0�@9�@UC�@L�@U�@^�@�g�@p�@z�?��|2HECKCON�FI� *?QG_Pv�1; L W_i_{_�_�_�_�_�CHKPAUS�1���3 ,�L�7�����ݿ�R?ٺ�:@"_D?[���\�/�_Bo ��/oioSo�owo�o�o �o�o�o�oA�[�O�1�?�; COLLECT_�2���t�4�wE�N K52�rbqND�E�s!�w�6�123456�7890�wL�pL��L
 H�/L)@�e��,?�Q��� (o����򏽏Ϗ�:� ��)���M�_�q�ʟ �������ݟ��Z� %�7�I���m�������-�t�2"�{ ��@�2�u�rIO #$�y�q�J6h��z�����6�TRP%E��p91�S�6�bq_MOR�3&v�< �L 0C4�C Ŝ��.��R�@�v�d���3��'��b/I?�A�A���L K��*L TP�r)�Ma�-�?�1�C߂�

�u�w��ܮ@x�6dߖ��`���PDB�p+jԥ�CPMI���� ��!� :�  3�1ິ5����J�\�'�V2��q0pq0q9��ߜ�g�������F���h��*0 �0 ��G��.���� �L ���mfdbg6�y�9z{�٠�UD1: RS�CH!n����DEF� *.xP�)u�d1:cpe�buf.txt��������_L64FIX ,��(���v� c����� �8J)n�_�������6H_/E -Q�</�N/`/r/�/�/@MC&��2.Q(�d�%�#��2/�-��45��/�?C:�B:�s��C��DC~��B�G�F�`�C@�50a�s�G� ��E��E�LJ��E�"5#]0�A=J����G�5+H��a�MƮ�G��2��0��n�  َ?��21�DT��P�4~P�q*P�ϴ�]�xNB&1�!`�B�V@|�D>��s�D!`Da�@��VfE��@q@Em��3J��E� E��3F7@E���fE��f�:T�>�33 ;�����@Gn�1��@o�5!� Q��f¦�A��T=L��<#�ޱ�Y���O��*RSMOFST (����2)T1�D* 2����2�
�A�q;��B�O�G?��ߚ<�M.TEKST��0_�sR�r!3l�_6�A@�j;@ �1�ACz04;@2�#cC��b��nR�p:d�
��QI�s4�]�QT�_��PROG ����R%.�o�T>�NUSER��r�a�q��dKEY_TBL�  .u�a|p���	�
�� !�"#$%&'()�*+,-./�w:�;<=>?@AB�C��GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������oq���͓���������������������������������耇��������������������
�i`LCK�l�U�d�`�STAT��S_AUTO_DO `���V-�INDT_ENB��0/�?P8�f*�T2v��eSFNc�5�]��GROU��6�-��Q%2����C��A��A��0���aa��B��=���H�{���D�@ �I�.��HE�W�i��{�������ß��STsOP[�m�SXC��� 27�jb�8
�SONY XC-�56�_�Q�����@�9�( А{�HR50����<�N�7`�r�ACff~��oԯ� ¯ ����A�S�.�w��� d����������п��+���TRLk`LE�TE�� f�T_�POPр疽b�eT�_QUICKMEyN柇�SCRE����i�kc�sc�ĳa�����RWc_��U�M���U 18Q <�܃o3���<�q� ��N�t߭߄ߖ��ߺ� ������(�a�8�J� ��n������������Cus Me�nu Edit �%custoy�n.stm��z��V�����v����� ��������A* wN`����� ��+a8J�p�����P�ounce Da�t/@ %GMP�NCDTA�L �'/]/�F/�/j/|/ �/�/�/�/?�/�/G? ?0?}?T?f?�?�?�?��?�?�?�?1OO��_?MANUAL��m�ZCDOb9IY�b�W�)TsW�O�O?|(��wCGRҀ:I[� B��$DB;COT�RIGW���DBG_ERRL&q`;֋�a�OL_�^_p_ �ANUMWLIM���`d�U�H`DBPXWOR/K 1<�[;_�_��_�_oo�mDBT;B_L� =��5���B4��@TADB_A�WAYS�aGC;P R=�עRpb�_AL�P��lb�BY��Y�Ph�n`P 1�>�K ,��\��'��F�n'1i_�MS�IS�{k@��@uONTIMV�M�T�bv�i
����fMOTNEND��h�{RECORDw 1D�� �0�CG�O��q�&� {b$�6�H�Z��xb��� ����я������� +���O���s������� D�͟<��`��'�9� K���o�ޟ�����ɯ ۯ�\����5���Y� k�}�������"���F� ����1Ϡ�U�ĿN� 违ϯ�����B�������-ߜ���/d�v���Ϛ߅����?�A�[��	���?�*�8�u��Ե�v����.����������I  �IJ�\���	�������%��������lbTOLERENCNtsB��b�`L���@�CSS_CNST�CY 2E([ a�arUeUb� �b������� /ASew������UDEV�ICE 2F([ ~*1/C/U/g/ y/�/�/�/�/�/1V�HNDGD G�(]Cz�kULS 2H-�/U?g?�y?�?�?�?�?�/WPARAM I�K�,'.%URBT [2K,8p<#/��` C��_ �v@�B�{`���CbATd�9ICut�Fv�0Ć`�F�rDyGKA��G����pd@�@�<�MIC��vW@� hD�  U�ĴpF�QAKH�K�XI ^qJU¾�c�M ��H�_d_v_�_�_�_ �_�_�_�_Aoo*owo�AC͵@D0C��G`�a 	 �B5�A��}�A��7A`��AW��Aݤ=��a�F #P�b�@�a�C>�<�aG B��BC�MB�S^�BT�B��2-�o�o�oHP��d� ��f fe� �pNv�=3CUo go�Oo}���� ���H��1�C�U� g�y�Ə������ӏ� ��	��-�z�Q�c��� =sڟ�ן���4� �X�C�|���i���� ֯��������B�� +�=���a�s������� ��Ϳ߿�>��'�t� K�]Ϫρϓϥ���m� ��:�L�7�p�[ߔ� ߸ߓ����ϱ߻��� ��H��1�~�U�g�y� ����������2�	� �-�?�Q�c������� ��������.��R= va������ ����<��%7I [m������ ��/!/n/E/W/�/ {/�/�/�/�/�/"?�/ ?X?j?��?y?�?�? �?�?�?O�?0O9? K?xOOOaO�O�O�O�O �O�O�O,___b_9_ K_]_�_�_�_�_�_�_ o�_�_o^o5oGo�o O�o�o�o�o�o�o 6!ZlGOuo�o� �������	� �h�?�Q���u����� ����Ϗ���R�)� ;�M�_�q���ПK�� ߟ�*��N�9�r�]� �������ß��ǯٯ &����\�3�E�W�i� {���ڿ��ÿ���� ��/�Aώ�e�w��� �ϭϿ�߇�0��T� ?�Qߊ�u߮ߙ�������$DCSS_S�LAVE L��������_4D  ����CFG �M�+���d�MC:\��L%04d.CSV����ā�  ���A V��CH��z����pm������  �p�����������y�IE�.���2�R�C_OUT N�!���] _ a�}�2�_FSI ?}� &� p������������ 4/AS|w�� ����+ TOas���� ���/,/'/9/K/ t/o/�/�/�/�/�/�/ ?�/?#?L?G?Y?k? �?�?�?�?�?�?�?�? $OO1OCOlOgOyO�O �O�O�O�O�O�O	__ D_?_Q_c_�_�_�_�_ �_�_�_�_oo)o;o do_oqo�o�o�o�o�o �o�o<7I[ ������� ��!�3�\�W�i�{� ������Ï����� 4�/�A�S�|�w����� ğ��џ����+� T�O�a�s��������� �߯��,�'�9�K� t�o���������ɿۿ ����#�L�G�Y�k� �Ϗϡϳ��������� $��1�C�l�g�yߋ� �߯���������	�� D�?�Q�c����� ����������)�;� d�_�q����������� ����<7I[ ������� !3\Wi{ �������/ 4///A/S/|/w/�/�/ �/�/�/�/???+? T?O?a?s?�?�?�?�? �?�?�?O,O'O9OKO tOoO�O�O�O�O�O�O _�O_#_L_G_Y_k_ �_�_�_�_�_�_�_�_ $oo1oCologoyo�o �o�o�o�o�o�o	 D?Qc���� ������)�;� d�_�q���������ˏ������$DCS�_C_FSO ?����-� P � �J�s�n��������� ȟڟ����"�K�F� X�j���������ۯ֯ ���#��0�B�k�f� x���������ҿ���� ��C�>�P�bϋφ� �Ϫ����������� (�:�c�^�p߂߫ߦ� �������� ��;�6� H�Z��~������� ������ �2�[�V� h�z������������� ��
3.@R{v|��C_RPI*�<������ �)��e���SL�@Z��/ 	//-/V/Q/c/u/�/ �/�/�/�/�/�/?.? )?;?M?v?q?�?�?�? �?�?�?OOO%ONO IO[OmO�O�O�O�O�O �O�O�O&_!_3_E_n_ i_{_�_�_�_�_�_�_ �_ooFoAoSoeo�o �o�o�o�o�o�o�o +=fas�� ��G����� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹���߹PIOC 2]OK  ��� )�;�M�_�q���� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������/ /+/=/O/a/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O��O�O��OCNUM�  �p��������RE_CHK �Q�{��A ��,8�rf_x_�Y 	 8b_�_�_���_�_�_�_o,o 
oPobo@o�o�ovo�o �o�o�o�o: Jp�_�_��Z� ���$��H�Z�8� ~���n���Ə��֏�� ڏ�2�D�"�h�z�� ����R�ԟ�ğ
�� ��,�R�0�b���f�x� ��Я������*�<� �`�r�P��������� ޿������J�\� :πϒ�p϶��Ϧ��� ����"�4��X�j�H� �ߠߺ���������� ���B�T�2�x��h� ������������,� 
�<�b�@�r������� ��������:L *p�`���� ���$Zl J�������� /�2/D/"/T/z/X/ �/�/�/�/�/�/�/? .??R?d?B?�?�?x? �?�?��?O�?O<O O,OrO�ObO�O�O�O �O�O�O_&__J_\_ :_�_�_p_�_�_�?�_ �_o�_4oFo$ojo|o Zo�o�o�o�o�o�o �oBT2d�h �������_,� >��b�t�R������� Ώ��������&�L� *�<�����r���ʟ�� � ��$�6�؟Z�l� J�|�������د��ȯ � ���D�V�4�z��� j���¿������� .�п>�d�B�TϚϬ� ������������<� N�,�r߄�bߨߺߘ� ������ �&���\� n���������� �����4�F�$�j�|� Z��������������� 0J�Tf�� z����� >NtRd�� ����/(/BL/ ^/ /�/�/r/�/�/�/ �/ ?�/�/6?H?&?l? ~?\?�?�?�?�?�?�? O O�?DOVO8/bO�O .O|O�O�O�O�O
_�O ._@__d_v_T_�_�_ �_�_�_�_oo�_(o NohO:o�o�o8o�o�o �o�o�o&8\ nL������ ��� �F�X�ro|� ��0���ď�����؏ �0��@�f�D�v��� z���ҟ����� >�P�.�t���h����� ^�̯�Я�(��� ^�p�N�������ʿܿ �� ���6�H�&�l� ~Ϙ��ϴ�VϤ����� �� �2��V�h�Fߌ� ��|����߲���
��� .�@��P�v��b�� ��`��������*�� N�`�>�����t����� ������8( n�^������ �" FX6h �l�����/ �0/B/ /f/x/V/�/ �/��/�/�/�/?�/ *?P?.?@?�?�?v?�? �?�?�?O�?(O:OO ^OpONO�O�O�/�O�O ~O�O_$__H_Z_8_ ~_�_n_�_�_�_�_�_ �_ o2ooVohoFoxo��o�k�$DCS_�SGN R�E��`��v1*�16-APR-2�2 08:21 �  <�Z��`2�-FEB-19 �12:18�`	p�	r S	D��NLX�qL�l��sH1NLZe�+qLMK�q�a��D׿W���~;
;;
�cV�ERSION ��jV3.5�.14	r�s�`EF�LOGIC 1S��E� / 	��w�@�y��@�~�rPROG_�ENB  �t��sp�sULSE � �u�u�r_A�CCLIM����s�!�WRS�TJNT��a��dEMO�|q�q�r�f�INIT T��z�J`�OPT_�SL ?	�Fx�
� 	R575��s̀74щ6҈7V҇50��1��2҄�x ��w��TO  E���xo��|V���DEX�d�b	p���PATH A��jA\1504�2022\R01�\ SѓPOIS�\ ӑѓҐ_V2�\ _�Ғ�{HC�P_CLNTID� ?rv�s �x�u+��rIAG_�GRP 2Y�E� (�r	 F� �F,D E�  E(p��D��A�v��B�  ����B����B���ά��C�eEC�  C�kI$CG�SCEZXB�GmA��f̐ 6789012345��q��@� ����=�A�V��v:�	qB8�y���� �u�� ��:��o߿�Fr��� �F���N��пj������*�<�N�A_��AZffAUG��AO�
AJ=q�AD��A>�R+A8��2��,��q��@�  A�`ApX�Ѧ�A�����`����G�
��`���A[��V{A�P��K
=AE��A?33A8���A2�\A+ׁ
	��-�?�Q�c؅�������xz�AqAj��c��A\Q�AT��L�וߧ߹��� ��c׭ϓ�yσ����� e���#��3�Y��� i�?�����������s� �B<�=���~�
����=�G�Q>8Qy�]��8��by�7�Ŭ���@�;�\��p����p@J�Ah7�v��<�C�<��
�=�w=����=���=��w2��;� <#���'��?+ƨCݖ�`(�Ur 4����I� U��A@	r?��� �����C�/��/=//a/s/	?�Tz�&�%���R �/G���R��%v��$��x��4E�4��
��J=CG�{CEY���.-�4b?P<>���3�1`�5��=�?�.ED��w�� �1D���3��0��S�<O���N��T	�T(UkT�]F󊆘��a?w������>�����W���ﶱ��1@����ڿw��E��BrLwDr�R�"Ao�Z3kO�/�A���AℲ�Bo3JA�"�OA\BF}OgB�O��B|IMI�3����g�c���� eO
_U8'__$_]_H_��_N�CT_CON�FIG Z`�|z�teg�u�S�STBF_TTS�
�y�Sip�q��ZMAUH���rM_SW_CF�P[`��  N��zN_��L��P 3\�y P; D?�E_a%�kl�g�k��?�3�o �o�o {�o�o�o (:#VhzH�8��|dPEN�� ��&�8�J�\�n�������a���̏���'"� ����6�H�Z�|d쏆���f���Ο@����P�(�|c]A��S�e�3�������#I ʯܯ��$�6�|dTILR�d�v�D��� ����п���ϐ�*� <�
��rτϖϨϺ���|fMUT�����`��2�D�V�|e@r� �ߖ�dߺ�������� �&�8�J�\�n�����R�Y���������1�|fpN�`�r� @��������������POMM,> bt������QG]�	�-?Q|fm�_���|eVAR�// �>/P/b/t/�/�/�/�PLI-��/�/�/	? ?-???Q?c?u?�?�?��?�?�?�?�?KEXO(O:OO^OpO�O �O�O�O�O�P���O _�O(_:_L_|f�Pj_�|_�_\_�_�_�_|dRE�_oo�_9oKo]o oo�o�o�o[��o�o�o �o#5GYk��IFY���|�����
�$�6� �Z�l�~�������ƏP�ޏ���Џ&�8� J��ed�v���V�����П��:b!� ����>�2�D�V��؇�p'v��������;���̯ޯ����"���}?B�T�����$DOCVIE�WER ]������	� ��frs:�/GMWIZMA�N.pdf UU�@�<CPUI�230_LN��   k��PlǴ $���ܟ���148_�I���3,	�� À/�oρϓ� �Ϸ����]����� (�:�L���p߂ߔߦ� ����Y��� ��$�6� H�Z���~������ ��g���� �2�D�V� ��z������������� u�
.@Rd����RC_CFG �^ĵ�!���������7���SB�L_FAULT �_�
J�NLTTBL 1`]�
 (  ac�4 not on ;m蒓���� �//;/&/_/J/h/ n/�/�/�/�/�/?�,�NGPMSK  ��e|TDIA�G aķϲ�j�JUD�1: 6789012345r2If1�*�P ?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O	?�G�e3�I��?_xTORECPK?]:
k4 ]_�7v[�?�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�O�O_�vUMP_OP�TIO��]rT�R�03a<uPM�ESF:tY_TE�MP� È�3B��K�p�A�pztU�NA�15�q=6YN_?BRK bĹ>2�yED_SIZEN/2' �ex�t�TAT�s�~EMG�DI�rfx�q�uNCv�1cĻ ��o(c�V���
��d�o�� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�IuN�`� r�����������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � Ϛ�G�Q�c�uχ� ���Ͻ��������� )�;�M�_�q߃ߕߧ� ����������%�?� I�[�m��ϣ���� �������!�3�E�W� i�{������������� ��7�%Sew ������� +=Oas�� �����/// AK/]/o/%/��/�/ �/�/�/�/?#?5?G? Y?k?}?�?�?�?�?�? �?�?O'/9/COUOgO yO�/�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�_�_�_oo 1O;oMo_oqo�O�o�o �o�o�o�o%7 I[m���� ����)o3�E�W� i��ou�����ÏՏ� ����/�A�S�e�w� ��������џ���� !��=�O�a�{����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����+�5�G� Y�kυ��ϡϳ����� ������1�C�U�g� yߋߝ߯��������� q�#�-�?�Q�c�}χ� ������������ )�;�M�_�q������� ���������%7 I[u����� ���!3EW i{������ �///A/S/mc/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?//'O 9OKOOw/�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_OOo1oCoUooO yo�o�o�o�o�o�o�o 	-?Qcu� ������o� )�;�M�goq������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ���!�3�E�_� Q�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�W�i�sυϗ� �ϻ���������'� 9�K�]�o߁ߓߥ߷� ��������#�5�G� a�k�}�������� ������1�C�U�g� y�����������M��� 	-?Y�cu� ������ );M_q��� �����//%/7/ Q[/m//�/�/�/�/ �/�/�/?!?3?E?W? i?{?�?�?�?�?�?� �?OO/OI/?OeOwO �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�?�?oo'o �_SO]ooo�o�o�o�o �o�o�o�o#5G Yk}�����_ �_���1�KoU�g� y���������ӏ��� 	��-�?�Q�c�u��� ������ϟ���� )�C�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ �����!�;�-�W� i�{ύϟϱ������� ����/�A�S�e�w� �ߛ߭߿�ٿ����� �3�E�O�a�s��� �����������'� 9�K�]�o��������� ��������#=�G Yk}����� ��1CUg y���)���� 	//5?/Q/c/u/�/ �/�/�/�/�/�/?? )?;?M?_?q?�?�?�? �?��?�?OO-/7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_{_�_�_�_�?�_�_ �_o%OoAoSoeowo �o�o�o�o�o�o�o +=Oas�����_ �$ENE�TMODE 1d�&e� + �P�P�p�q��Q�u�U�r�xRRO�R_PROG �%�z%�VE�R� �TABLE  �z�,  �@ ��] ? �  ���� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ� �ϻ���������#�� �SEV_NUM� �r  ���q , �_A�UTO_ENB � �u�s�_NONZ� e�{�qD�_  *������%������P�+�ж�8����v�HISA��Q��po�_ALM 1]f�{ ��T���P+��W�i�{��������_OUT_�PUT 2g�����P2�_:�|�  ��{���r.��pT�CP_VER �!�z!=���$EX�TLOG_REQ����mـ�SIZ\��{�STK������}�TOL  ��QDz���A= {�_BWD���d���_DI�� h&eo��t�Q<�STEP%7|�pQ OP_DO����qFACTORY�_TUN��d�	D�R_GRP 1i�yj�d 	)���p�� �[����N�#.T�&hB�( ����-�>� C+<~B��_�B�7�B]�]B���Bu�ICB>6`B� ,�BPiA�|��A�M�Awa��k8|`>�A��woA��Aӣ�A�e�\A�A���M���i��m���ˠ��ejW��T���6��S<���>C&`M'�R
 �GE{�{K%A�N���.�������/�/�/I��=N�%B�ƈ5Co@UUU'?UU�/�P?�/ E�� �E�@z3x1�4CO�HcGP�2L��uS�1K�y
�C?B�\?L����2�18Q�?&{ffC:G:��5�9{���5?>F�? <>��6��I��E���U�I�9�:� EATURE j&e� �Sp�otTool+ �cH oduc�English �Dictiona�rylA�R��4D Stan�dardeH R5�3Analo�g I/OdIMI�G �Agle S�hifteHII)��Auto Sof�tware Up�date  av�ad�Cmatic BackupjI�Qground EditinglA�
IF�@Came�ra�@FdIVLO�A8Pell�Lm@�
EN8PnrRn�dImShER69�18Pommon calib U5P�kBdcol�Vsh�WQgF04 R�\cyo�@lAt\j7�W��@pane�S F� O�Xty�@se�lec�@ OAD�7Qon*Q�PMon�itorgYons~�@t Path^�ntrol Re�liab�@kBlf{va�QrnerY`�g a�W04D�ata Acqu�isckBuct\~�`iagnosQ��AiDENDI�as~^bFaultshE�fd -�bpen�se Plug-�i�d4SDocum=e<`Viewr`jC��P5�`ual C�heck Saf7ety�Q (�@tA�hanced M�irr)`Imag�e �@"0xRob� ServY`q ovcro0xT1#`�dad704�`2vUsr`Fr;P�Q�`t@�xt. DIO V`fi�d `p�rWend8pE=rL�b� mPD�x�ws  I.�`�sr�@�p ���eVIFFCT�N Menu pv�ac�VFTP In��pfac��@,p�G#Pp Mas_k Exc4pg�q��CHT/�Prox�y Svt�Afr�d�igh-Spe�8pSkizT�!�d��`�pmmuni�cP7`m@g����u1r��pdILo�A�A^2�conna2lAwPar�pInc@p�8`r�`�fdjog�KAREL �Cmd. LY�u�Dp�v�Run-T�i�pEnvlA" �#�PK�p�P+Ps�	PS/WlAjui?.Lic�br�v
! k`�pBo�ok(Syste�m)�EEq�@MA�CROs,��/O�ffseaRIN�T��H grip�pr`c�SlAWel�@MMR#`b�hQP��pMat.H�@l�-QOp�c "MF��PMechStoepj�t`��wm~�L;t�K rp@$�x8px�@	PfGPCVL��>wqSwitcBf9�#iop֔�a.�p�TOfronx���m��8pC֔k�filvY��Ox��@g ie�n_�M�`i ApCpl8�^a*a;�n�`
�E�`p�b�T�rꢣ-TQ�-SjCD5RP?CM fun��ߣnk_�Po�dr,� ORDEX�ua��}r�a 88 J<�Kri<`FC�C�A�>k�g NumZpa�xc XPʡ���p �Adju��iE "x[�ʵ�J \ars@�tatu�fȣʵ.^ABoxiD_�ȷ�yR��`RDMVqo}t}@scove�AN�tRem��qn�G�  y�Z�[qc�_qu�est ������o�pxuF�X@N�PX bP�eNSc�hedule0 �(S=0) ct3rl6���Seq�iDp<�X@�BLibr�CjC�`��C�@:uP Ц@�X@om�t�ssag,��tZA�jD�xB� �C��hEclP<�Ӈ�PredC��B�/I0� .pc~��TMILIB��<ȣ/�Firm�BfG�82.��P�Acac$P,VX���TX^Z8�S�`��eln����O0
P��_@ ���gFt�@h�r�� S�imula(aAQ )9d�h�ug�P�VbdCcs��#P_a��&���v. 5��U�SB port �PiP�p;a sl�ds��nexce�pt8pt�a�  H�59���xfGs\s��PVC�Qr��� ER H,�`8��Gcus�`J� � q���PJ�SP CSU�I �4c?���XC|�Fp�Web�a�e��rs�`��[q 5Pˠ��r�2t�a�p�`����_\���Gri=d_�play�t��X��T��iR/�.�J�oDR-2000i?B/100P/�����@Graphic<���ADV-��?bAC���h���� �p��Alarm C�ause/r�ed|�BlSAsciij��ͲЁr`d
Upl�р
ؠ��DQ�@'Pxai�AOT�B�sRec��k��QQ�2�ere6p CkW�O�rĊ��ccsu_�CRT/�Keybo�AMaQnDpC^bH���Ag:�Coly@ aG�u�F�t�PPƥC�yc�@4���orix%p:�e�DCS Z��./����!g2.Av<#!q�B߅'�c�P�DH�cJ��DRAM���A(`���	�g1s1�;��a 2&P�H�A���DP�`N�q[q.�cTVSP�s���Outpu�B VcAR�qd�D$M�!therNet��!tm@TYLs�:2Q�OSnif��tBR9&B2ca�*` �A�RA>`�p�����@� ��p8qs��@D���uG�RS Cհomi�z5�t���2�Ͱ��P�M��adi���<PAk/R���3Z2y�/�2X9�*�8�#1��M� ��p5q�i�pxmyp���Util2"�@�rNRT:N"P�COn���l>zX    �@���5�ݐb�����PCL1�&�mh<��0CX��vvB��1<�FA_�Pay.Id�`�"x�$2U߀f�Б�P����FLtr�u��k�cZ���qا��k�d�peq A�pymP���R
�<8�&ROS V6!�e�cSN/�Cl��t�c��[pi�pN�o?V�ģ�Jump����o0�F.	�����PEED OU�TPUT�/��!/FILE�&�d�rR��s�u�Zero �Down'#��i�R�)ص 64MBp�b;�<�bFRO�k�X/�lb!�� p�u"#t�d?TW�>&s\H#� g1�D���!Q�+�Ds�x�tr�l��nT p0MAI�L���FE� ��[ pS@C�r9ցAdp�0d�V5�ts0ݰ�!H��M G4 GMP�ucٴ��IABIC\��ڳmpmwL�@�ar7l �Ec�MaIx����eQ��BSH ξcro���PH7WAY�� g �W�~��RS4�?'�g�mp� Ѝ�p�!yn?.(RSS)C���ires x)_�ZÈ �O{�S�`�]��SuS�@e2tex�8��W�KaLimRw���l������S��P�OpQ��c SWI�MEST f��F� 00Y��@��� �"����>��9�Z� �U�/��q����� �� ��K�=ů�X��ru���\r�:�ysh.4����@Q��y�����≿���mwiz��Ƴ�0@����S���E�5���a�g�.�D�0�R���sLϺ�|�h���� �ϦÌ��ϟ�& ���� �B����a`���1A� /�A���e�3߉����� ��ѯ������+�J�sszpE�f�ra��zp��}��t���[��wr�ϙ���pt_ ���	�*�g�$� F��A�W��]�w�� y���,R���U���W� q���S�Q��ﳝQ ԺP!���=���� ?���)���`sQ� |`�r�` "�" ���8Z	�vAp #��"��g^�p��sre/ϩ�.v�isv/�,�wi P/R�d�v���/,φ� �/��<�?`Ϻ�L?�� pςϔ��? �?6 HOl~HO������O��O�O� #1O/E�rs+OE�QJVO! syD_fS-}�d`_�D0�/�Uad"���_#II)�_�Tmp?Y�n"Po���!/?�őAo# H�6\o~c6��xo~%6pۿE%�_Ϸ793�oNF$ H7�o�d1�o��h#oBt22�o�g3<;zt3 H8t�s�825�ET "<��s, Pa��st\sl�f�O�O�XF -�Qo�oao��litk/�_#��5�G� �c?�73 9(�:�) "_)���r�fd~O��ex	 ��Rߙ�#5&;�X"���!���xeK?R��pC�}%H�`h��Ol�~�|&- k���?o�����ngl$��}�u�?UVc�ї�FLX��"�֯f|&Pa'_�5cf� ��+o��Ҕt�TW�h�e���gVtFI�){��l&_������~spÏUUD@�$�ZDin�/ɿۿc1tK��c�Trc�E%�3.�Ж����
�XPL��TC�5�!<��6�U������TX�/}%"SG����J64�o5�t�����uif8��v�Pri�/=�nd��}%�g����6eT��i��� ��~$4���4*2<u��}%SeG�5f3EN�$.f��=O�����os���� �WG�oϤ����#arO�S�W��@6��2&his��u$��H/��zdG/Y/�..3vrO��u51��`�����Vrt�/ ���D?f3 k��/�>E .�?��=} �?�?`N� +/9_C� s[�2p�y�GP��DSvgC?e=�;��O�  ��Ach`�OퟷO!o��ta�_fQ�uc/��CVg�]�?r.S�ѕq�?� o nce_�GT�8oZcmir_vdc�t\+�!�l`�o�EbK�800�o�o(_�:_uBUz?|tc$�ep�_�Fg�߀�3RI�_i�ra��y������s#1"O@e9t�O�67\k6�B�P\0�
�uO��V�Ȁfo��aZ�(�\f	_���fj؏�O��_M��_~hu�?�'!p�/�7�O�5b V���>��.pc��Ecf/Evc�o�_�)�<�?�� cmo_���<д���Co���NToo�5on�q�F�x��Ob�fd -\�f��F ����R8W_��5RC���ί�gf�#��ӿ�w�  �H590 � 990\\�21~�R782b��� \�5a�j748�J614��H�ENATUP�V�q L��545�  ��R��6���VCAMV��CLIO:�����R�I�� ����UIF.�� IIt�6��]0s�CMSC�Ј����� "Ms�STYL  ��|��c28���p��636����NRE*�\im"��5������3m��nt�SCHFaw���DSB~��PLG��brDOCVܲ#|�CSUVAr7���9!��P��ORS)Rr���8a�c蠌��0���EIO���BC Jt�54y� J8Же��q.��SET�F����/Basi��7����MASK���PRXYR��7n�`\et\�OC��CE"����-���;���fcb��б�f� "�����J53�9R�HW�\cW�L[CH�CC:�Os�rD�0-�P�MHG��Mg]�PSt��Ms҆T�MCр���D�T:�D�D�MDSWڢ�D4�at^�OPd4��R��T�63)�[pp�EN
 P:�361)�D�60a�P�PCM��ms^�Ra0H�h�� �50)�t+��Щ�S:�=�5�0��L�RS��gd2Z�5��j�69)�T��FRD��|�RMC�1�IW:�S��D�H{93I�SNBA�`�alW�[�a���SLeC��\P��HLi�7_cm��SM ���Nе�PPu�_f�n��2	N ��H�TC��_ma��T�MIЁ�At�q�tl p PA��_r��TPTXj�TEL 1��`���q�c� ���8x��t�m�H���9�5!�w� �)���VUEC�\�� �FR� ��H�VsCO��T�VIP�9c� ��SUI��$�X��r�WE%B��i dT��	��
��2��9�d��GzLsDIG(��lPGS.�IRQC���w�6x�l��t�6��d�t�8��bh���`��g�66����7�Ѱw�t�8�6m��J9\�7�i�@�)�<�l���Q�s��AB�nt�p.��3��J68���P�2-�nd!J�56(6!�#R5"Xh����1m��8 �!@/J75��8N )�D�6��@� �B�q�� �v���BАa��Щ�t����7���76a��)��#R5�8N�y�D��gJ77m��57)�v�54)�dmmg!̳"T69���$64Jm�s�$5y��1y���� q��$87!6N3VD�Ь#R7�X����EQ��!�! �h��R6��F-2A0��Xᐱ@2-�9386��a����y��3H�����7�04!��\h82�D�F2eBK�7���D0��fdRFWB5.f�_BS�� Ctl��TO��r����wORD��DLP���840'�7�1Lo�a_JNN!�(F��NN)��@. !ћPa�54a��GsMP���IAB)nch3�N�-�l�N�`����q�n pf@�PHpA,F�� �y<(�)�   �"��j��CPR�0p� "�p�6D10�6~�ETS}ka�reM�� KAd�°/�p CP9м���Gene�R�I=��� �UREL�Vmp,�V䱤U�\=�ldp\�UT�RAN�UPy=�t�\ka�Udpcp��U�q�_�[`��UqPl�@g��=�-��=�Gu��@=�͠�V:!�U45� H�VH�g863ޯV7 H7�UH7+79�f2�i7�f�@t�V�`6�f811�U�68�h�0�UAIC��hR8�V80�f"�@�f (C�Vx`�V��A=���=�90�gE��U8=�sfmn Hv$�xvq��e4~�=��j693fhSw�xb�3&g�@i�U(�Patl� TXP�f�)esw�$i ��p�v! jwOB�VJOG�U�B�U��t=���J��Mac�U@�AfJ�	�U��uo�  �U�=��"=�_耤UpxfBPert.�U/F  !Xh�U���Ume�VH�R Jn#vH62#v24�j�#v855�V3�i6�42�f�x�`0�f3U8�V6��0v4���f780�Vp�i#v�7	��d�g1�` w3�;v!��i;����g68�f5͛�f0���b�w19��h�v79�gh�D��
w1��Иw2^�
�h2�f2�`И�f'@�שk�75˧��w�1�1#�k��f4�k�0(Ʒ����3v35��f�62֧й�_Z�cl�b�oriC�II)ػVX"��23�VMN!SӆPBM�&g3iAY�GCur�VI�[�Jʧ�MPof73 ( �oas�v @����X�o���X�NT^�v9vone{fng�_,m\pRw�pK� �a��д�4�u���f �p�ϖ@�д��Ќ�E�:Y�h]�01SS�8��(��V15S�_
a,�0IuPOvX `d��p�x�P���tet8ۖ�r�t053��.�����P�ߗ�18��Џb�cse�v�1�a���8943�l 	U�v�0RL���	@��ail�V �d�JtR�LUH�P@X�i@K�7��L�uJ ����LVW�nĀHv�����ߔ\mp���57��Arcw�2�e�1Me	A9�R f�@C��5���\h�� "T8[�( �obt_��"�	rd8�2F����40��5�fq�#vS�erv�Vk2�DE%R�VIPЀ�5;v�@���V�B��s�intz�@�j&'hq.f���89�V����\�sWf1�s�ltkxL��@9� tkr�H/Z�gtpfQ@�V0]@?� �Vntj��z�7F�M-wace,X�)��p�;v��j89�fn�h?6�\mtfHi����4�oWf	 �:  H59�@��`A�21Z�v��@8I2G`A5eD���P�1%Q��anA�TUP�
�@5�45�dT�B67�VCAUP,��CLIO'�@RI��D��@UIFNdsKhi�@6�E�@I�@�MSCN�0R�D8��STYL2� v�A28Z�B/1 Q;63�JNREJw Q]5�D-50R3uD����@SCH�'�@D�SB��5PPPLG~6�DOCVj��p�PCSU.�0i�A Q9eT�`FOORSRN� Q8eD�H804�A0�U3��QEIO5T�р@5�4�DlC`�D5XB]"@`SET�p�P�J5�Ep70�PJ�7�EA/1�PMA�SK�tR H�PRXYf$�`R7���QHOC�D�S�` uT�S�@�D��7�beD��SJ6�E�SJ53�9�YHv��R�LCH�d��`�VPW-70�A0uT ��F�`HGEd�Ѱ`S�UA0��`�V81�`CDUdH��b0�D�cJ5�U:��D�`DSWJ��q�e (P-Pq�e<!�qR�D�ѠR�d�`_pMAEN��B�dH�d0beD \p�`CMT��1�@0D����b�D685�s�dā�b�D��\�b�d0m\r0�Dp�@PRSudPa�eU��B9�d���FRD�DE �@RM�C%�g�PPf15L,`@93u(PPNBA��^q�PeD��PPLC�D70l.FPPHL�T��PPMd�pc�P�DcSPPUtH71�b2eD Ѡ�ܥDSHTC�Dph3�@TMIUT�B�%t�TPAEdC-�fl�TX�ITEAL%��Sbp%t��e�@�8�Et�BuD��@9�5eTAC"�A95��}rUEC�dc "?PUFR�Dl!�A�T�0\c�PVCO4du X�@IPUT���@SUI������X�Ed�SWEB�D}�3r��T�D�CR62�D7\c4��CG��,��IGĥL�2 �PGSF�IRCUT`�`@�6��"CSL�A6��u �qR8�u�9p��� we��rP���\�7del�R��92�ΑR86uDg I/P���<�ĵ�C�P�d�SMa"p��TAB6��se�Q53�D,�7J68�Ej9/���6�dTX^�56e�R�eTprsmPa�Sܢ�eTmke�`R7�1uD��5dU\sm�k�a5��,Ѡ��d23\s�Ad�(A���d =�P%t<S�@���@@�v�CR`��\e7�e}BJ76eDL�r��d�cmp_�R5T�縢��RUd\ik���77uD��R57.�d83\�r4�d����j78�―���64uD�@�`�PUdԣ81Uj��%ts=�8�7eTL�NVDudt�y^�7T�|sFREQ��<���eTm��dvsj6�4uPEE�p ���d����dm�?��@�Ud94 (���DTPU?�$���"PeT�@v�R8�UNTSo`�b���M�D0d�tc�s�PF���CBS8�Tm�/`CTO�D	 `�@�PEd��QLP�T�CP S`��ion?�NNU墐p��d�� �eT��4eD���@wGMPudredPgIABŤ�T63�j,�P�Dpp�qS� 6��PH$�L�"P�DRS���rP�2��p�@P]RE�g R?pRS�rfaA6�խPoasTS5�L�SLMud�f=�6$�L�Ð�Te܌ ��ene�$rs�1}$x�s^��t�par�	 A�	4<���g AW�	� t�	���	\��<R�awaw 2fTET�
\sep��VUR]�m��s�ch�-�L`rcMs�	FL�`p/d"/VUN�O,sh`/dr/�H�/lp/*̼/.+TO�/`mo�n ??VUC�, A�RC0*�<\?.+62D.;�0O�	- _*E͡��9ݡata�
�e�tJ����)p\a�	�±?��]`J��B�\b�9�OJ��N �	̂�܂�Irn��9���847�:Mq�����	<��K�*3B7.?�
b7�Zܒ8���M-4�
������31���9P<�lM1\m4���h6�:31"�	!e ~khs�p:/3�
Z� H@joa�[1�pi��OcXM_j���\pfmPj��_#_��_����500,pz-�1y�`�ZM����0 "�j��/ZL<�/Z42�k�]6�8�	Sec�
�o~ �j,>Pb�f|�`k�PR�:H.�a�, \�
�=825�J#< ��O�X���_*hs_f0*l�0� �*�`�:�ok48.kTR,/Z�=h���:\���,�"�
r� ��3V_, �o\�i�{iA/_�D� x�Z�`�	-100�
# I����A�h���I�сj\_*<�63.x��܀/Z10F/���RDϊTlP�	(R-�jTUD��{�j���{s���20Xޫܟk25.kF-�"�:7M�_�q�7�j��v� p�j0iBo����ά25/�}�|Pȯj����5���	 ���@�bY�{\߾�30i�|����P�:제@O�xph�?A�4!3o�ݼ\��
6܀�J�A�66ߊingN/ZA/2�
loh_�U�?Jnu����.��-43ߪ
-�����8/ZS)��j|�0��ߤ�_��� �Esth�\�793��&�ierO:�)�_��ui�V�d\g/J��� cy�le x�Z�ߊ22 S�zM�R5�Im�����tpcy ��:t\dN[m��\�etn��=��4 H J�9�J77_Z75�9/Z85 �6 �R��J9ߪJ87��zP3M2+S� R_[S0O]�z9;90�8 J��m-�R8R8��l�6�03/Z�J,�Ki�pe?��si_�P����gs�ZLMip�NlMip�[���t�egOJ\�89�+8�4�+� 9�Z����(�In  �STD��m�aLANG��dE�qdEpfpmdE��F���dE0\fpdELS�E�FR J5dE!� PrdE��F! �TdE
ELS�F"�C�Flly dEJ�760dEated�dE�dE�dEt\j�7dEc "F�FP�CVdEL�dEmc.�v�F��dE|dE��dÈP0V�HV�bsw�GNDdE5�5.fdEh754��FMawV4S
�dE��dEM�V H7��Fte 2�FPa �F��l_� ���WzOhA�flr�W�O�S\t�bTV̀�_��SVLR; Mf/7LdE�ѐ<VL�dE��HdE�Pe��Fm�dE"��_� r7ldE���F�dE���Kv3ܰdE��dE75;3\dE.pc�f�i��dE- L�F0i�D/�O
�Pf���GM�adE/7H,dE)3 "�oI�\l�FܱXf-��V6\�x6gf0�1dv�P�vh.�F�Y�� Wv�dE,�i�WI�_V758�͠/V �(�LR-`�r�LR4vD[�g�vh_fC�sw.�N,�vfd��87�W���pRB}T�EOPTN�tx���r��-350��Aaक|�����h�� "M7�������N��74mӖ��E���h68������M-�71�����H64��Lo��49 (��50E,�����A��9\m��8�핐<�4���-�`��0AHV�b��bY�5��iC/�\���0Ӗ{h6Ɨ75H"������̰��Ф��PIxܦ|���670.�'0iCĨw�H����l�ܦ (ۧWS���0G�D��0\��R yq���r�����,��}�W�1�����DPNh@\�\�7Uq]�Հi\��[�S$p\��xs�`r]�\gws�Ɛ�a�ŝ�^�1lph�"@g���\��\ŝ-\�/70W�Ǣ��Ů� ^ø�^�I�ǐ^�lC�ŀr`uŅA]�e�g�q�T�\żR��fgwr-P 6��������  ���R��ss�pc��! ��PC�:P�� ���R R6� �593��44 =R�� J78���P1 �� �81�m��T���nter`��8R����t\�׏mov.������ snl�P��pnl�ׄ��5q�a|�a(gistx��is��lsvw��a)��1o��8�J�in��b���30;���ge�n��p�a�H$�H52��8�������CH��A���v��)v*���B%�R
�%�m�a696z���or,���z�A#�H574�ռD�aadv\��A7DVS�IF�������	! aw0��1�$�In+����651��9�Qi ����A`� �4���fm�ٍPo0	D4`����H/�M@�845�����@b��0Ma�Y�41lf`�pr`��A4fm2�@�a%坡�����5���U-�4h( ��22aLg&d�� ��03�����!'��r�/� h���`w�Rm�ormP��M�Q/� m��C��@6鑝�21[���M�����1l�祱ADJ364��"\a��P�/�*2l7�R�ՙ�8���%�120L�t����C�`�5%q�1qM?�0iFTr���i�pfc64�?' 4?�,4\�7H?Ac�?�?�G Ov�a?�]  ����ݢ�� PT�698�9���YS�t M1e8/J/�&csc6�Iw skc7! j$�=T�'g. &0�7�95/�90��cD�CO�1 R/�R88c1�`X2��%!S6��%��d7R�����oub[�& Pxw����_ \j9cD_�n�z�]%A_C�tr��5��0	st�n?tioorIe��1Q1��G�5x�:��3�hH54�g]�]Owon gVe�O8O>�p�ZPH�֌�o�Vcse�d�op�tim��d\o#zp��܏�h?�y�nd��cm�� f1u�`��CM�g�`�������(w�p���,\���W�O;Sm\c6t���杠���p����Mw�kF96���R7k�81��56�hS06'70"�h 	pFp�F�T�i/{*etd�F���	����@_�E�'�	���j61�6gle���M��c�u�/�4���6j0�.�V�����!�Э��Ƹ��-W�JĬ� �L�I�M�?�sm�mai�[�PI JNN�99B����$�FEAT_ADD ?	���q��y�   	 ո�ϔϦϸ�������  ��$�6�H�Z�l�~߀�ߢߴ�������d�D�EMO jq�   ո+�!� 3�`�W�i������ ��������&��/�\� S�e������������� ����"+XOa �������� 'TK]�� ������// #/P/G/Y/�/}/�/�/ �/�/�/�/???L? C?U?�?y?�?�?�?�? �?�?O	OOHO?OQO ~OuO�O�O�O�O�O�O ___D_;_M_z_q_ �_�_�_�_�_�_
oo o@o7oIovomoo�o �o�o�o�o�o< 3Eri{��� �����8�/�A� n�e�w�������Ǐя �����4�+�=�j�a� s�������ß͟��� �0�'�9�f�]�o��� ������ɯ�����,� #�5�b�Y�k������� ��ſ����(��1� ^�U�gϔϋϝϷ��� ������$��-�Z�Q� cߐ߇ߙ߽߳����� �� ��)�V�M�_�� ������������ �%�R�I�[������ ����������! NEW�{��� ���JA S�w����� �///F/=/O/|/ s/�/�/�/�/�/�/? ??B?9?K?x?o?�? �?�?�?�?�?O�?O >O5OGOtOkO}O�O�O �O�O�O_�O_:_1_ C_p_g_y_�_�_�_�_ �_ o�_	o6o-o?olo couo�o�o�o�o�o�o �o2);h_q �������� .�%�7�d�[�m����� ����Ǐ����*�!� 3�`�W�i��������� ß����&��/�\� S�e����������� ���"��+�X�O�a� {����������߿� ��'�T�K�]�wρ� �ϥϷ��������� #�P�G�Y�s�}ߪߡ� �����������L� C�U�o�y������ �����	��H�?�Q� k�u������������� D;Mgq ������
 @7Icm�� ����/�/</ 3/E/_/i/�/�/�/�/ �/�/?�/?8?/?A? [?e?�?�?�?�?�?�? �?�?O4O+O=OWOaO �O�O�O�O�O�O�O�O _0_'_9_S_]_�_�_ �_�_�_�_�_�_�_,o #o5oOoYo�o}o�o�o �o�o�o�o�o(1 KU�y���� ���$��-�G�Q� ~�u����������� � ��)�C�M�z�q� ���������ݟ�� �%�?�I�v�m���� �����ٯ���!� ;�E�r�i�{������� ޿տ����7�A� n�e�wϤϛϭ����� �����3�=�j�a� sߠߗߩ�������� ��/�9�f�]�o�� ������������� +�5�b�Y�k������� ��������'1 ^Ug����� � �	#-ZQ c������� �//)/V/M/_/�/ �/�/�/�/�/�/�/? ?%?R?I?[?�??�? �?�?�?�?�?�?O!O NOEOWO�O{O�O�O�O �O�O�O�O__J_A_ S_�_w_�_�_�_�_�_|�_m  h %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �//+/=/O/a/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳�����������  �	�)�;�M�_� q����������� ��%�7�I�[�m�� �������������� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m�� ������Ǐُ���� !�3�E�W�i�{����� ��ß՟�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���'�9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}ߏ� �߳����������� 1�C�U�g�y���� ��������	��-�?� Q�c�u����������� ����);M_ q������� %7I[m �������/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�u���������Ϗ ����)�;�M�_� q���������˟ݟ� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻�����(�����
�-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���� �����)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	- ?Qcu���� ���);M _q������ �//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_��_�_oi�$FE�AT_DEMOIoN  d�E`��`-dINDE�X:kIa�-`IL�ECOMP k����{a�Hb(eq`SETUPo2 l{e�b?�  N �anc�_AP2BCK �1m{i  �)h�o�k%�o`~`Be�on�o �!��W�{� "��F��j�|���� /�ď֏e�������� +�T��x������=� ҟa������,���P� b�񟆯���9���� o����(�:�ɯ^�� ����#���G�ܿ�}� ϡ�6�ſC�l����� ϴ���U���y�� � ��D���h�z�	ߞ�-� ��Q����߇���@� R���v����;��� _������*���N��� [������7�����m� ��&8��\��� �!�E�i�t�i�`P�o 2�`�
SYSSPOTg.SV�*L�TEM*d� %���K�o/) �7/�EAL����/�&/�/J/\/n/�/?� /9?��LSCAH�/�/?�?� .? �?R?d?v?�?O(?AO�/�0IO�?�?O�O�!6O�OZOlO~O�O�%_0OI_�*.V�R ��_ %*� _�_��_�_cXP�Cp_oQFR6:��R$o1i�_Uo`[T�X�_�ogv`�o�ixDo�o�*.FnPzo%	c�a-9xq�o]�kSTM�o@�b`~q��yL��kH��w�4�p�X�j��fGIF� ���u����G�܏��fJPG����u
�<�0ˏ`�r�eVJSxo���� 4�S��M�
J�avaScrip9t͟��CSS�&��u�D�O�Cas�cading S�tyle She�etsQ�� AZ?*.BIN ��?FR5:\��̯�S�AutoZo�ne .bin �file}���DAT�������P�߯��dat���ARG?NAME.DO���p\��Z���̴ݿz��̰DISP�տ��: �`��R�a���
KVAREEGW�9�ǲ��b�\�	��POS��<�ö(�����ύߛ	REG\����ȱ��j�|� ����B���0��� �|���9TPLINd��� %ȱ��r�����TPEINS.XML$�L���:����%Custo�m Toolba�ry��9PASSW�ORD���FR�SVн�|�%Pa�ssword C�onfig���9WPAT�mQK[@�X� %BU:�Spot App� Proc z�a܁�gmc��.v����������Fp���� fg*��_%H`�%�Wiza����gmpncdtaN�Z��
Poun�ce D��GMWIZLO��/��pP/����Log"��at�m���%��/����tio?n GRS4?��MPBk?SX5p?�}� MHPLG�F>��?�?���?O8P��OCO�?gO �?xO�O,O�OPO�O�O �O_�O?_Q_�Ou__ �_(_�_�_^_�_�_o )o�_Mo�_qo�oo�o 6o�o�olo�o%�o [�o��D �h���3��W� i�������@���� v�����A�Џe�� ����*���N������ ���=�̟6�s�����&���ͯ\�� ��$�FILE_DGB�CK 1m������� ( �.�UMM?ARY.DG ��ݧMD:4�t��0�Diag Sum�maryu�"�COcNS�"l�O�D:������� sole� lo"8TPA'CCN�S�%;�x����TP Acc�% tinϦ�S�6�:IPKDMP.'ZIP����
����|����Excep51�߲�`�MEMCH�ECKn�տc���~ !Memory*/���ބ)o�RIPE�]�o����%�� Pac�ket�!	�Ӈ{B���ST^0���߼��
� % �S�tatu�<�	F@������t�	�����mment TB�D���e-�)ETHERNEV����C�T�����Et�hern)�ur�42��< ��DCSV�RF���������� verify� all�Ԧ�=X��DIFF�����0diff�QC���CHGD�1�y�  X�GRk��	28�� 6�ZGD3���(/� �O/�U�P�0ES.�?n��FRS:\l/�-��Up�0es L�ist�/��PSRBWLD.CM�/�p��"�/�/��PS�_ROBOWEL2��,��I��?/��?����Net/�IPJ a.����()�0GRAP?HICS4D�?�?��?�?%4D �Graphics� File����ch��SM��O!O��O��A/Emasil�?���r2NOTI���O�O<_���Notifiqc��`O�˅�r2?SHADOW6__�-_�_��Shad�ow Chang�_O���r2RCMERR�_�_�_Fo���`CFG E�rror Det|�@�_ �J�CMSGLIB>o%o7o�o���e��� xX@�o�`��)�`�ZD�O&�oJ���ZD+�ad�oyl���)<pIRDG?_REPOR��/|AS%iR���nour Repo}r�/ ~�DB�PRCSW�p����X��rSpot �App proc'ess��&���p��9�K�U}e%p��og ��?��MP� ���ȏ]��MH Plugint��	�Sh��&�	�>�<P�b� h%x����`VAR� ڟ�ԟ��d Varc{hg��basei�>m7TPDRA*�B�T��`u�� �x�� s�\)��A�x�x/�l�����Z� ������ĿS��w�� ϭ�B�ѿf���Ϝ� +�����a��υ�ߩ� �P���t�ߘߪ�9� ��]��߁ߓ�(��L� ^��߂���5���� k� ���$�6���Z����~��������$FoILE_� PR� �����������MDO?NLY 1m����� 
 ���_�VDAEXTP.�ZZZ��q�H��6%NO Ba/ck f]@ "�ͽlN��8��� �H�'�K]� ���F�j� /�5/�Y/�f/�/ /�/B/�/�/x/?�/ 1?C?�/g?�/�?�?,? �?P?�?t?�?O�??O �?cOuOO�O(O�O�O�^O�O�O_)_��VI�SBCK ���*.VD*_t_\aF�R:\CPION\�DATA\__����QVision VDu�_�O�_�__ o_Bo�_Soxoo�o +o�o�oao�o�o�o �oP�ot�A�9 �]���(��L� ^�������5�G�܏ k� ��͏6�ŏZ�� k������C�؟�y�����2���ӟh���M�R2_GRP 1�n���C4 w B�)�	 �������E�� E��@ڣء�s���O�HcGP��L��uS�K�y
��?B�\?L���+�(�8Q�?&{ff�:G:�O��9{��[��A��  w���BH��C���N��B�ƈ���s���ѿ⽬�@7UUU��UU���0ϫ�>x'>C��q>F�;��E�=���3� �9�{F:�4��9˽:N}��:LG:�%�Ϙ�[ϕ��Ϲ�������{�_CFG {o��T !��b�t߆�1[NO ���F196�839  /]RM_CHKTYP� B���)����������{OM��_MIN� �'���	���X���SSB8�p�� ��6�%�-��V�h���TP_DEOF_OW��%���>��IRCOM�Ў���$GENOVR/D_DO��
��THR�� d��d���_ENB�� ^��RAVC��q�VQ �ϥn�Y���}�������� ��!�OU��w���)������8�?���-^/  C�y >iX���"�AȑB� ��©�	o�"�SM�T(�x/���,�x��$HOSTC8�1�yL[�Z� 5	NNN#�~�e��� �/*�2/D/V/h/���/ 	anonymous�/�/�/�/�/? M_qN? �/�!/�?�?�?�?/ �?OO&O8O[?�/�/ �O�O�O�O�O?!?3? E?GO4_{?X_j_|_�_ �_�?�_�_�_�_o/_ eOwOTofoxo�o�o�O �O_�ooO_,> Pb�_s���� �o�9o�(�:�L�^� �o�o�o�o����  ��$�6�}Z�l�~� ����ŏ������  �2�y�����K����� �¯ԯ���
���.� @�R�d�����ϟ���� п���;�M�_�q�N� �����ϖϨϺ���� ����&�8�[ϑ��� �ߒߤ߶����!�3� E�G�4�{�X�j�|�� �������������� e�B�T�f�x����0�ENT 1z��� P!PLC � �����!�124.11.2�40.31���! �,��	G|? �c���� �Bf)�M� q���/�,/� P//%/�/I/�/m/�/ �/�/�/�/�/?L?? p?3?�?W?�?{?�?�? �?O�?6O�?ZOO~O�AOSO�OwAQUI�CC0�O�N��4��O�G�O!192.168.���/_�IR_3_�O�_�@R�outer�_4_!���!_uCPCJ�OG�_�_��IT�P0��O�CCAMPRT�Ho$o�PIV1DoUgR�TR�oto�o�o��N�AME !��!�ROBOao�oS_CFG 1y��� �A�uto-star�ted��FTP��q���G�� ������:�L�^� p����'���ʏ܏�  ���Xj|Y���� p�����şן����� �1�C�f��y����� ����ӯ�������R� ?���c�u�������r� Ͽ����:���M� _�qσϕϧ�� �� ��&��Z�7�I�[�m� 4ϑߣߵ�������~� ��!�3�E�W�i���� ������������� /�A��e�w������� ��R�����+= ���������� �����9K] o��&���� �FXj|~P/� �/�/�/�/�/��/? ?1?C?f/�/y?�?�? �?�?�?/,/>/�?R? ?O�/cOuO�O�O�Or? �O�O�O_(O)_�OM_�__q_�_�_)�`_ERR {z�_�V�PDUSIZ  �#P^T@��T>~�UWRD ?Fu�A�  guestV%o7o�Io[omoo�dSCD�MNGRP 2|�Fu�P�XA#P0��@�#P�#PK�d 	P01.03 8�1� �`M�0�  ��  �`l� pj�; ������������$���������(p�}  
H�Dp�Dp�  ?jDp�DpT��lp})lp&����lp�zlp�4��0�*�`~�`��c
@[r��+ p$p�$p/� s��b8{`�f�seL�[p{�\�d�o&�k_GWROU�`}�Y�`��b	�a�a1W�QUPD  �pC�UY\���TY;��]��PTTP_AU�TH 1~�[ �<!iPend�an�g�@_� �!KAREL�:*�
��KC�1�A�S�)�VISION SETf�����#Q'�ȟ���� &�����c�:�L��p���ЄCTRLG �]�u�u
#P��FFF9E�3��DFRS:�DEFAUL[{ � FANUC� Web Server����QӁo d����������ɿۿ��TWR_CONF�IG ��k �f��QIA_CHKCMB 2��g��Q ��!OROBO.�p����w�w�y@�����` �������b`p����(]��ρ�w�z�Ϥ� ������9��σ�B� '�#Q5�G�Y���}ߏ��߳���5�DEBU/G �C�
%�t���q�����(�D�EL �C���8�?S�T���1�ELB=�m�S�<� ����7�+�=����� ������������R
 .@�dv� ������* <N`r/��� ����//&/8/J/ \/n/�/�/�/�/�/�/ �/}??"?4?F?X?j?��?�?�?�?�?�?0�F�OBJ 2�C�᠊����ڑ  n��E`!RBȨG �E�A�OWN�s�D�O__�` 8�4�6�  6_X_Z_l_�_�_�_�_�_�
Pi�ck Press綋O�F�AŷHJm�O  _�O�o�oxo2_�_�o �_�o(R<^<�
kDropo~o �o����9�K�]� �o���v������Ə ��ڏ��&�lD��+� ������s������k� 5���+�U�?�Q����u�������U�2�GR�P 2�C���ʕ�����	 < *�L�~����������� �Կ��2��:�h� N�`Ϟψϖϸ����π�����R�<�i�0�'@�  ��v@������0���$f�� ��ѿ�?�z  Ć�C��ؿ�=aɔT����/  Ap���u����'A���� �Ԃ � 2�Ĵ����Ț����@@���f��������ؙ�|���� ��������)���\�Q���t�ZHN�p�r�:btJ߰���H��� �� N8Z��|�����
����B:6f  m�6 �?a3Cdq�`{�Q�ɕ�=lCLCFG ��[  3����O����_F?`i�i��,�k����m/*/ �OGw 2��
 l,/a�!PO�/�/�?�/b/ �/�/??'?�/9?]? o?�?�?:?�?�?�?�? �?�?O5OGOYOkOO }O�O�O�O�O~O�O_ _1_C_�OU_y_�_�_ �_V_�_�_�_	oo�_�-oQocouo��NET ����f�UM_CHK  ]_�c��f�ELB�o 
�fFOBJxD!5&woPAIRT �f�WTu%tOTF ���?u D/ � BH  =��c�A3�
�qr2��� ��t  t!k��'ӟ'�9�K�� o���R��V�h�ُ� ����!�3�����
�{� ����b�t�՟�J�\� ��/�A�S��(����� ���r�����ʯ+��=��o�SETUP ��H<���K��
 	
P� ��o�o�o����ҿ ��"�C��<�>�P�rϰ��a��ѕ������������2��O�X��=!����Fq2��_/�Q�
Z��Sp�� �;!+�$T��Z!C��"�	O�)
7�Z!O�]����V���������eO����6pa��i�"���-6"�Q< ������< V��="�< ���$�Sp�"� �$�:�����+�"��s"�< ?*��"�K���OKp"�c�R�R�a���}�?`�Epim"�B�V��"��#CԦ�^�)����"�%+�6p�p &,���`�"�'m�A�*"�(���"��d"���|����e��e�"�+�2��"��@���#�5��G�U� l��x �ϭσ��Ϗ������� ����7;m Wi��k���� �!B7iSu �������/ �/S/2/O/q/s/}/ �/�/�/�/?(?�/? O?9?[?�?;/u?�?�? �?�?O�?O9O#O5O oOYOcO�O�O�O�O�O �?�O�O5__A_k_�_ __�_�_�_�_�_�_�_ o	o+oUovo������� �bWTPR ;3��{
 ��o}��~Э��d���o����"�dc��b]�x����x��2"s�o�o�o �"4FXj| �;������� �ˏB�T�f�x����� ����m������,� >�P�b���������� Ο��򟟯�(�:�L� ^�p�����A���ʯܯ � ��$�6��Z�l� ~�������ƿs������ �2˧`B_CHKCMB 2��i�4�dek�ROBO�T��G͸� 2�y ��RżŒ�W�b��V�P�kߕ�(�2�z9� K�]�o�j��%ߎ��� V���� ��$�6�H��Z�l���DEBUG ���
���+��Q�S�:�w�����L ���M�Ooqoso��ELB��Y����� ���������v� 3EWi{��� ���x�A Sew��,/�� ��//�/=/O/a/ s/�/�/(?�/�/�/�/ ??�?9?K?]?o?�? �?$O�?�?�?�?�?O��O5OGOYOkO}O��F�OBJ 2�����1�P�HW���no�E`��B�OW MUYQp_�N�CJT�_�_�_�` 8������ Mo�_'oo3o]oGoio��o��
Pick? Press��2_DVYQ�^X�mm_�_�_ BT�_�o�o� ������/��kDrop�o%7�� ���������wA� +��7�a�K�m����� ��͟�l�p�ҏ3�E� W��,������ܟƯ ��ү�����2��.��@�R�����GRP ;2���Ee�8������	 <ѿ� %�[�-�[�A�Sϑ�{� �ϫ��Ͽ������� E�/�=�_ߍ�sߕ��� �߻����� 0i��@��  �v5@�BÝ���CQ���F:� �Eᰥ�z  ĆSS�ᰤDQ�p�TE���  �ApS�����A�vE�� W�  ��Ĵ��i��u��fZP@��C�¾c� �Bv�@�#�5�v�Y����}��������������g�������ARt ��W��ߕ��� ��+L#Esp]��
��eR:6f  ��[ ��a�Cd�@��`R  STYLE103_TC��$���p��MSHAN�D 2���
��0�c���/��y/�/ �/�/�/�/�/&?	?J?���G�n/@?�?�?�? �?�?�?�?�?-OO"O X?j?|?NO�O�O�O�O �O_�O�O;__0_fO xOJ_\_�_�_�_�_�_ o�_oIo,oKot_�_ XojoLo�o�o�o�o! (:{�o�of xZ����/�� $�6�H�����t��� h�Ə����=� �?� D�V���������ߟv� ԟ���
��.�o�R� d������������ #���*�<�}�`�r� ��ſ̯����޿�1� �3�8�Jϋ�nπ϶��ȿQ"LCFG m�]+  ���A������3�d�<#�,��5��[��"O� V��`�9���OG 2M�], ld�b�!� ������4�����	� -�?�Q�c�
�u��� ����v�����)�;� ��M�q�������N��� ������%I[ m&����� ��!3EW�i����F-NET ���� 8��?����Q"PA�IR 2�]+ �������� P��Wҵ�x/�/�/ _/�/�/�+C/�/�/(? :?L??p?�?�/�/Y? �?�?�?�?�?$O6O�? �?O~O�O�OeOwO�O �OMO_O�O2_D_V__�z_�_/��SETUoP �������s�KP
 �	
ڰ&��//�� �_oo(oJoxo^o�o@�o�o�o�o�or�Y�v��+��0Bz}2~  �P��Q  �PFTNђ�_~t��ZP5G�B��w�zp�$P���t�r�	R�x
�t���]+Ь��Z���t�x��xЌ�t��aZ+І���+�6r�Qx��q)�"�x�V9�=r�x��J�XЙp�r�B�`��X�:b�^�Z��zpR�sr�x�?*Pr���FpmpKpr�������a�p�̆{�O�imr�R����rб#�t���p)�Բr�%zp�/r�&�+�K��r�'�p���*r�(P�r��dr�	�|:�1�e+�e�r�+np�p�r�.�@���r�������� lxpx �o�oҟ�oޟ�)��� �P�:�\���h����� �����ܯ���:�� F�p���d�������Ŀ ����� �B�l� "�\ϢρϞ������� �� �
�,�V�w�J�l� �߈ߪ��ߊ������ �(�R�4�V��r�� ����������<� ��,�N���n������� ��������8< nXz��^_�e��iR �WTPR ;3��
 ���QnR�p�E%{RRkQd��"��lQQc�W2q);� _q������ �///%/7/I/[/m/ ?�/�/�/�/�/�/�/ ?�?3?E?W?i?{?�? �?�?^O�?�?�?OO /OAO�OeOwO�O�O�O �O�O�O�___+_=_ O_a_s_�_2o�_�_�_ �_�_oo�o9oKo]o�oo�k� C_3D_�CFG ���O���b+r�AZ_CALIB� 3�9{������}, ����/�A�(��e�L����������f?ROBOTʏ܏ �|���X���|� c�������֟����� �0��T��N�r��� �4�¯H���H�� � =�O�6�s�Z���~��� Ϳ��񿀯��9ϰ� ү`�毓�濷Ϟ��� �������5��.�k� Rߏ�ϳ߮���N�p� rτ�r߄�U�<�y�`� r��������	��� -���:�L�������� "��d�������; M4qX���� Z��x���(I�� ��x���� �/�3//,/i/� v/�/8�/�/^L/ ?/??S?:?w?^?p? �?�?�?�?�?O�/O =O�/�/dO�O�/�?�O �O�O�O�O_�O_K_ 2_o_V_�_�_4O�_�_ ROtOo#o�O�_Yo@o Ro�ovo�o�o�o�o�o �o1C�_Py�_ o�&o�&��� -��Q�8�u���n��� ��Ϗ^ʏ���� >��q�ď��|���˟ ���֟����I�0� m���������,�N�ܯ b��b�3��W�>�P� ��t��������ο� ��/�*�S�ʯ�� � � ��ϸ�������+� �O�6�s߅�lߩ�8� ����V�h�zόϞό� ��o�V��z����� �����#�
�G���T� }�������<�*��� ��1UgN� r����t������$IC_AZ�_CONF �����FS����� ��k�<��7MEMB�R 3�F HROBOT������� �$///B/l/N/`/ �/�/�/�/�/�/�/�/ ?D?&?8?b?�?n?�? �?�?�?�?�?O�?O :OdOFOXO�O�O�O�O �O�O�O�O_<__0_ Z_�_f_x_�_�_�_�_�5PROG 3�F o�_oVo ho�o�o�o�o�o�o�o �o%.[Rd� �������!���*�W�5SCHE�D 3�F  HR������d��
�_��XVoxel ?Sched1��������ƅ2Ϗ�:���!3�)�����4_�q��ʟ��5�������6��Z���77�I���B��8���꯽�9ǯ(ٯ2�bÉ0�"� {�F�Ά`�r���Ɔ� ����̿Ɔ^���� Ɔ��8�J�\�Ɔ� �Ϥ�Ɔ6�������Ɔ ~��"�4�ƆƦX�j� |�Ɔ��߲����W� ��J�9��]�� �����/���"���w� �j�5���Y���}�� ������O���B�߀1�U��y���3 '���o�	b-��l�PACE 3�+k ��_�[�T� 	 �YD��  E	� D�e��B���C��� �P,�P  �?aG��F��_ L/����/ /�/ D/V/h/z/�/�/�/�/ �/�/�?�??.?@?R? d?v?�?�?�?iO�?�? �?OO*O<O�O�OrO �O�O�O�O�O_�O_ �_&_8_J_\_n_�_�_ <o2o�_�_�_�_o"o doFoXo|o�o�o�o �o�o��o0B Tfx���X�� ����,��P�b� t���������Ώ��� ����(�:�L�^�p��� ˟����u�ܟ� �� $�6�H���~����� ��Ưد����˿2� D�V�h�z�����Hύ�LST 3��4 B�ػZ�@ϟ������� �����b�A�Sߘ� w߉��߭߿������� ��+�=�O�a�s�� ����������6���'�l�K�]�����f�D�P_CONF ѡ�JP
Wd h��ؾ��E�Ez���;� ?8Q�@7��ͽ��`�I���SCHED 3���
�D�eadlock Prevent�� 8������� ���E8 R{n����� �///./</e/X/ r/�/�/�/�/�/�/? �/?=?0?J?s?f?�? �?�?�?�?�?��hz �?=O0OJOsOfO�O�O �O�O�O�O_�O_&_ 4_]_P_j_�_�_�_�_ �_�_�_�_o5o(oBo ko^oxo�o�o�o�o�o �o�o ,UHb ��?O�|��� ��(�Q�D�^���z� ������ʏ�� �� �M�H�R���~����� ��ݟП��� �I� <�V��r�������¯ �ޯ���3���� {�n�������տпڿ ���.�<�e�X�r� �ώϨ���������� �=�0�J�s�f߀ߖ� ������������&� 4�]�P�j������ <�N����#��0�Y� L�f������������� ����$UPZ �������� (QD^�z ������ // /M/H/q/����P/�/ �/�/�/�/???6? D?m?`?z?�?�?�?�? �?�?OOOEO8ORO {OnO�O�O�O�O�O�O ___._<_e_X_r_ �_�_�_�_�_�_oz/ �/�/�_aoTono�o�o �o�o�o�o�o& ,]Xb���� ����#��0�Y� L�f�������ŏ��ҏ �����$�U�P�Z� ������"o4o���� �� �>�L�u�h��� �������ԯ��
� $�M�@�Z���v����� ��ݿؿ����6� D�m�`�zϣϖϰ��� �������E߸�ʟ ܟ6ߟߒ߬������� ����.�4�e�`�j� ������������ +��8�a�T�n����� ����������& ,]Xb���� ��`�r�#�(F T}p����� ��//,/U/H/b/ �/~/�/�/�/�/�/�/ ?? ?>?L?u?h?�? �?�?�?�?�?�?O
O�$OMO@OZO�O��$�IC_DP_SI�D 3������A� � �OwF�O�O_ �O_<_3_E_r_i_{_ �_�_�_�_�_o�_o 8o/oAonoeowo�o�o �o�o�o�o�o4+ =jas���� ����0�'�9�f� ]�o���������ɏ�� ���,�#�5�b�Y�k� ��������ş���� (��1�^�U�g����� ����������$�� -�Z�Q�c�}������� ����� ��)�V� M�_�yσϰϧϹ��� ������%�R�I�[� u�߬ߣߵ������� ��!�N�E�W�q�{� ������������ �J�A�S�m�w����� ��������F =Ois���� ��B9K eo������ /�/>/5/G/a/k/ �/�/�/�/�/�/?�/ ?:?1?C?]?g?�?�? �?�?�?�? O�?	O6O -O?OYOcO�O�O�O�O �O�O�O�O_2_)_;_ U___�_�_�_�_�_�_ �_�_o.o%o7oQo[o �oo�o�o�o�o�o�o �o*!3MW�{ �������&� �/�I�S���w����� ��������"��+� E�O�|�s��������� �ߟ���'�A�K��x�o����$IC_�DP_ZID 3ߥ������ d �� �������(�U� L�^�x���������� ܿ���$�Q�H�Z� t�~ϫϢϴ������� �� �M�D�V�p�z� �ߞ߰��������
� �I�@�R�l�v��� �����������E� <�N�h�r��������� ����A8J dn������ �=4F`j ������/� /9/0/B/\/f/�/�/ �/�/�/�/�/�/?5? ,?>?X?b?�?�?�?�? �?�?�?�?O1O(O:O TO^O�O�O�O�O�O�O �O�O _-_$_6_P_Z_��_~_��DL_CP�U_PCT�P�QB��  �P A5;.(�SMIN�\��� >�c���GN�R_IOERR � �S����ICD_BG ����U�-iicmedCbg�_Sochdd�X�4gi?o�ocl�toiisv>o�obo��o�a�o3�o:`o �o�oXjq"�F~�y)ud1:�����bDEF 1���|a/b-�q:`��pbuf.txt����a_BND_BOX 3���;-a 8����XΏB���CF`�#m�b�V ���P �D�V�h��X
3�����Wd��|d�ub��Z�STATE 3�.�� �|b�����(��L�;�p��W ^�����ï���֯��X��;�*�_�N���r����X��׿ƿ��@���CϏ�b�#o�����~���O�АSI�`�j�yh�TNPT^��M_DOff�" �ՐL_SCR�Nf �e �T�PMODNTOL�.�jE�_PRTY���Q^�VISg�E�NB.�� �_F_FRCVRm���<^֧�M  ��3���Ϥ�RSMPRG���������$IO�LNK 1�� ?�~����������b�MASTE`���eOSLAVE� ��_�_AU�TO��	�<�UOPxJ�@�E�YCLEk��;�8�_ASG 1������������ ��(:L^p�����Y��NU�Mc�
=�IP�CH��|�RTRYG_CN�Pb�O)�O_UPDc}��e1 =�h��������w���PP_MEMBERS 2����` $ԇ������ԋ�#�PR�CA_ACC 3����  T�v�  ��� 	��@ -� 7ߕ��P5�P&�&?b� }r#/$�
2_�RD,�BUF001 3����= o u1 ޕ o u0� 0o�@�$`�#p tX� � p�$p�$p`�u:K
*0p���$��$��$��#q�� �_@q u�<td �q� 7� >q�$q�$q*�$q�$q�$r� 02�$r�$r�$r�u�1]�Xr�$r��u;2�BLr��$s� 3�AXs��$s@uC,�H�xs`uBbj��s� 2�B�s��u?u?  s��uCt� �s��u>u>�  u�@th �t uBI�+�t@�#Ut�$t�$t�$t�$Ut�$u54u�$u�$�u�$u�u< A�T�u�u6��VAu�u6i�m�u�$v54vl�  l�n�$Un�$n�$n�$n�$%n�$n�$s)2�/�/��/�/O &�!Z{
�" pT��! �A�!�B� �A�!�B� u<�@??)?;?�@t� �T1�A\1�Ad1u;cP�Dt1yR�@LyR�0uC�0�0u��`�1yR�8�R�8u@�  �0�Q�1�A�1�A�1�R��D�1�R� `h��?�@��A�B@	QAu6�@%@)b�D 4A9b=@>ADOVOhOzK3�O�E  �C�`�B �`�B�@�B�@�d�#�@ � �b�"�@�"�C�b�" �Cr� r�dS�@�d %S�@�d5ScPtEScP �dL3cPU0Br�dd1Br �dt1�r�d�1�r�0�r �d�1�r�0�r�0���1 �r�0�r�2�S�r�d�3 �S�r�d�S�@�dC�@ �dA�@�%@��d 4CCc��McK`�d]cK` �dmcK`�d}c2���;3��� 4�į�����qȄqҮ�HIS}"���� �! 202?2-04-11�� }�=�"��� �(��b"�8��< �P 9� H   1� j�L��@� ) !`�h��p   & &  2 ����<����T��`�J!��R� b� 6� -�?� ; ��PP�]���j� �- �@ 7 �
u�P�}� : ����x��; ��J��  	���?@|������*������u�"�T�ߚ�����	�����������@ , M����P��]��� j����@��u���}��������i���q�1_�P(y���?@2��R�������9W�]��&��?T��D���4{�U��  4T�ߚ)3ɯ��I 	�K�}�@
 3 ����/���V=� .΀Ly�,�?@��e� `���������������]3��TT�ߚ2�|���,  I娟 % (���2T�@��M�7K�Z�]� _�@4�-�?�/- NU�<���u�c���T�ߚ�b�'��	I �@P��_�j��p����%��"�T�$/  :E֊ߚ�b a�s��K�H��rJ�]�@H�j�H��bJ�u� }� H�i�H�M�H�y�H�Q� J����������@��৿ݯ����� !� -]�'  @JA�8g�[�@`�QQ��+���"  7 ��u������ϟ���p�R�d�%A�=(�Pl�]�6ƀYA�l�S�@0)�O�����i��M���y�p�	 ?@aX��S�Aں� K�9o������F� ���߰����╿ ���e�l�"4F Xj|��E�r��$�p�^e���^����`/ &�"./?�_�Q�V/h/z/C�U�C�`� �/���/��)/?M!�.� `2?D?V<	Aa !�3�E�W�i�{��� �����������`�l&�`I2[hTUhT hT(hT0hT�8 2]kQ@�TH��TP�TX�T`�Thz�Tp�Tv 2_kQ ���_oo]Z��nQ yqvQNbPNb�PNb�P Nb�Po@�R�q�Q�q�QEE�TI�T�b�PK�T�OkQx 2�A�� 2SkQ� 2V�kQ�hT�hT�hT�jhT�hT�hT�`iSl�`I-~kS-�sS�-�{S.-�S.g��S.y�S.��S.m�S/#�S/\�S�/��S/��S0z�S0~bx 0w�c�0��c0��c1��c1G�c1}�c1���c1Rr� 1���c1��b�aH)U�kS)jr� �(; )�R0 )}��P�)Q�P)٣S*��S*J�S*��S*-��S*��S+�A�`�+a�c+��c+���c+��c,.�c,lu��`,��c,��c=->��`-C�b�/�aH%kS%ZQvP%d�A~P%�A�P%��S�%��S%ۛS&z�S&�bP &��S�&��S&��S&���S'�`'o�c'm��c'��c(
�c�(B�c(z�c(���c(��c(��c)Q�bs?aH 6������ ��(  �֋S!�S!~b@ I!�A�P!
Q�P!�r�X "�` "Nz�S""�p "��c["��c#$�c#�Ro� #��c#��c�$�r� $?�c$� $��c$�@�bOO����Ε6�0��U8��@��H��P��UX��`��h��p��Ux�����������U������������͸���`���I_�CFG 3�:[� H
Cycl�e Time!a�BusJqd�Idlz���mi�nk��Up|v�|�Read��Dow����
@���q�Count>|�	Num q�����k�!`���S�DT_ISOLCW  :Y�� m>G�_USED�PV��t�J23_DSP�_ENj�����OBPROC��rB�����G_GROUP� 1�V��Ad8�?�Bg�ψoV�e0�=�!`Q S�xߊߜ�[����������ge�o���IN�_AUT�`rB��P�OSRE�ώ�KANJI_MAS�`��Ċ�KARELMON �:[(�!by��������
��h���W��:Uİ�d>�Y��KCwL_L4�NUM�W�z�EYLOGGIN�p?P�����F��LANGUAGE� :U����DEFAULT� ��(QLDX��@L��ī���>���G��I���!c���PU@� �!`']G�  �?�,��MC:\RSC�H\00jq����N�_DISP ���Ϋ�R�P�&OCT�OL� !aDr�^�A���GBOOK +���d!`��662�BVhz ����������		� ��/���_BUFFw 1�V� �qb,ʅa/1\�}/�� �/�/�/�/�/??? D?;?M?z?q?�?�?�?��?�?�?
O���DC�S ��� =��zq�	\N:UrO�O��O�O!DIO 2��� ?P�O?P@���O�O__)_9_K_ ]_q_�_�_�_�_�_�_ �_oo#o5oIoYoko�}o�o�EER_ITMS�d��o�o  2DVhz��� ����
��.�@�8R���bSEV|���M�fTYנU��oຏ̏ޏa�U�RST���ESCRN_F�L 2��M@�� ROR�d�v����������TP��Sϩ�N��
NGNAM�ī���n�UPS� GI��r���-�_LO{AD��G %�%PRT50���1_Vt%��$M_AINT_V�?\�?  (%��į �в��֯���3�� W�B�{���x�����տ ������/��S�>� w�bϛφϿϪ����� ����=�(�a�L߅� �߂߻ߦ�������� '��K�]�H��l�� �����������#���G���XUALRMX��;� 炅�b�3���8�;�A���C� ��I���0�����_GRP 2]ƭ� �q&	���"9�  } ��l$A,>wPH e����� � $HZ=~i� ������ /2/ /V/A/z/]/o/�/�/ �/�/�/
?�/.??R? 5?G?�?s?�?�?�?�? �?O�?*OOO`OKO �OoO�O�O�O�O�O_ �O�O8_#_\_G_�_�_ u_�_�_�_�_�_o�_ 4ooXojoMo�oyo�o���D_LDXDI�SA��0���EM�O_AP�E ?}�
 ��k  2DVhz����FRQ_CFG� �����?�V�@�4�@4�<��Cd%�|��~������4� �16-APR-�22 10:12�:24 2�>�6:�02R�H�27:1y0n�H�45:3���5B�00:04:28�������0�� ��%��o.����:�L��^�T�Q�T�R�T�SeT�U_�T� ����V��,(HOME_?IO 1 Cl�-� ���ڟ����M�4� F�X�j������Я�����ۯ�*�]�ISCw 1��k �b� m���u���9�������5�C_MSTR� ��k�SCD 1��m�ؿR�Կ v�aϚυϾϩϻ��� ����<�'�`�K�p� �߁ߺߥ�������� &��#�\�G��k�� �����������"�� F�1�j�U���y����� ��������0@ fQ�u���� ���,P;t _��������//:/%/^/��MKƵq���qp/$M�LTARM�r�:%��" [#*���/�$�`METPU��`�s���NDS?P_CMNT�%�p>� ��N>�#��qf?p45POSC�F7�&�6RPM�?�9STOL 1���k 4�r#�
�1Y!�5�?G�?O 
OO^O@ORO�OvO�O �O�O�O _�O�O6__�*_l_VQ1SING_CHK  ?�$MODA�s��/��)�YDEV� 	�j	MC�:���RHSIZE��m�ȦUTASK� %�j%$12�3456789 �GoYe�WTRIG 1�K�l����oz�0�o�oz�)fYPaz����SEM_IN�F 1�%�`�)AT&FV0�E0�oR}):qE�0V1&A3&B�1&D2&S0&�C1S0=A})GATZR��tH� �aq�o��xA�*� �N�5�r��� 8�� \n����'�^� K�]����<������� ۟�����ď֏�Y� d����Ɵ��n�x�� �����1�C���g�� ,�>�P���t����� �ί?���c�u�\ϙ� L�^��ς������)� ܿM߄�q�,�6ϧ�b� �߲�����%����� ����2ߣ������ ������3��W�s.�ONITOR70G� ?�[   	?EXEC1U#��U2��3��4��5��Tj`��7��8��9U#��`����� ��������@������2U22$202<U2H2T2`2lU2x333����QR_GRP_S�V 1�'{ (�^Q��X"����?����`������6+l�1a_D��n�!�PL_NAME �!�%��!�R-2000iB�/100P, B�ase �}$RR�2 1����0�|0	X d[/�//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?G?Y?k�2��?�?�?�?��?�?�?OO+O�R< x?UOgOyO�O�O�O�O��O�O�O	__-_�PDDOU^
D_y_�TPh_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �_�_�o�o1C Ugy����� ���o�o-�?�Q�c� u���������Ϗ�����)�;�M� �E@ D�  �Fv�]W:  �z���aRdv�^��� ����ߟ�_�R�k�ד�$�5��X�[�  H�s�i�{�������ϯ��:���$������`�^� M�W� �@D�  k�?��q�W�?aPs�aQ@T�;gk�_T���;��	l��	 �� X�X��5������, �,�X ��:K���K��eK��ɜK~o�K{�GK�M:�ࡿt�3�=�:?���?��S�@�
�_��%��I���`���;g=�X���X�����������  �ô��l����  ��w*=��@�N���o�H��π҄��G���*���h  �� � �WЏW����c�G���$�	'�� � ��I�� �  ���;�:�È��È�=�����'�@������]��j�]�!֔*�8�r�N�m�O  '��:@���?�6@���@X�@����[���B��  C����B�l���6\Ӑ�B����
 � ����e��d�H�!�B����'�k�0����D�aQDz@�f� �ϊ�u������߭��������  ��� :]��  �,aP�?�ff��!3�� ��gy(�����
�ѳ"�(aP�P����˳˴�5�ϲ;���;aʤ;�D��;��;�	�<$D�@^�QA��,郲]�?��@�?fffs?&�}�A��@�,�,���x�� �s��q��a��R '//K/6/o/Z/�/~/��/�/�/�/,�F 0��/)?�/M?�n?�X@?�?<8E�0	��vf�E�0�E��2 �?�?;?O�?8O#O\O GOYO�O}O�O�JJ��M�O	_d?*_�8H^��Eƞ�G���~ƌ��ĳ�׽���C{�O�v_�_�_�_K��IZ�����_o�_P0ooTo�A0�Al� wb���Q�o^�Ho�oDg >��@o�o�oz[���Á-D��?D�` Ca*Z���p�q�q����W~COLCC���Ck�B��1B-v�=��������)���1�W
�u��^�����
��7
=AX��Blz��X���������ic��ö�=BU(���f����LI��JJOޔLU�W�H�� I%�K�A���M�DLs�L]���HP� H�R��k�U���8L�iPJ�
`H����H���A� �����ˏ��(�� L�7�p�[�m�����ʟ ���ٟ���"�H�3� l�W���{�����دï կ���2��V�A�z� e�������Կ����� ��@�+�=�v�aϚ� �Ͼϩ��������� <�'�`�K߄�oߨߓ�`���������Gj�,���D��{4����Ā�RZ�a�CB�߾�������_9�����C������F��r(�q�`������{�3��1�V�0m���q3Z�qb�������v�������v3�g����!�;�%?D93ҵ�	�[Im���eP;P��A�O�Q� 
4XC�^e�������� 8�`t��"//F/1/�j/�O�/�/�/�+�-�/�/?�/;O��?)?  �e 3�C??�?y?�?�?��?�:  2 EiMsG�"�Fvx`��tB�ata�`C@D
��A�p@�oIO�pE���rEј F���vC�> G� �GED Gt$ ?F� E�f�_O�O�f�?O�O__<&_�s?�ff?Q�D*�1�d�p�pb!9�d�k
 -_�_ �_�_�_�_�_�_o o�2oDoVohozo!��b�����0���$�MR_CABLE� 2ݿ ��tT� b&
�o �	{)�`��c1� ��Cy�as�� ����-���?� u���]�o���Ϗ���� �ۏ)����;�q���Y�k����o�����ڟ<�N�`��*��** �cO�M ��i�}��� &+ ��g�%% 2345678901��Bҥ �������j8A��
��}1980/�0B� 00:J� �*��W��TESTFECS7ALGv�eg�J8Aid���
���� ��b������̿޿� 9UD1:\�maintena�nces.xml��-�   
��`	��DEFAU�LT{(�bGRP �2ᤪ \ wym�6&��� �1st� mechani�cal chec-k�����@�����5l��J����x'�8ݎ�H�р���controll#er�Ͽ����ȱ�`7����߭�G�M���"���'�.��5������y��|��Kѻ CX��2���J�\��0��B����Grea�se bal�r bush��������������X����Cc�V�oling fan������������j�C��ge��.u�t/teryj3Y��!�@���5	fx�:L^��$ e�gp�{(f���!�!��5,�� //t9��
caKbl��@W!<�`_!f/�5
���/�/ �/(/:��W��
W/?]3�/�/V?h?z?�/�:�Overha�u� ��2 !x�`�1�?��6?H? 
OO.O:�DOOBO �k�8�OkOɕ�O�O�O WO�O�O�O�O_'_u_ �_c__m_�_A_S_�_ �_)o;oo�_!o[o�_ o}o�o�o�o�oso�o �o�o1C���c�HIST 2�ꅕ�p���L���c����jJ�K�5��5� -937.�2 hours _RUN 9]��u W��(�:�x��p��_�����I�"�L�hYn�-3227.6��������������qo���������p"��S�e���q����=�tI�N&Y�N��908��a�p��_�����Ӄ�wP�hI��6768.4���p>/�P"�����DR�hb��87	5��`�
Ę�,v������e�SKCFMA�P  �uN�p }����>�ONREL��`��	�~��EXC/FENB;�
���T�FNC[�M�JO�GOVLIM{�d��s���KE��}�z����_PAN:��²���:���ûSFSPDTYP{�F��SIG��=��T1MOT��J���_CE_GRP� 1�u	�\$�	��ϩϐ����9 ���ϴ�!����W�� {ߍ�D߱�h����ߞ� ����A���e�w�^� ��R����������+��O��8�PD_�THRSHD  �$�F@ f�QZ_EDI� }����sTCOM_CF/G 1���~�������� 
��_AR�C_X�����T_MN_MODE{���f�UAP_C�PLj�NOCH�ECK ?�� � ��� ����,>�Pbt���{NO_WAIT_L7����l�NUM_RSPACE�����/�$�$ODRDS�P:�f�OFFS?ET_CAR��[�J&DISW/H"PE?N_FILEv }�����)!PTION�_IO��ʱ� M_�PRG %�%�$*�/�.�#WOR�K �|�i� ��p)5�;� v $�C0�M4A��8C1�xA��* R�G_DSBL  ��w	���?�xORIENTTO:�f|�C���A H"�UT_SIM_DR�'��"* V. ?LCT ��$����d+LI!@_P�EX7 y/?DRAT�7 dUMO UP ��O
 �p��O�O�O�O�I�$P�ARAM2u�����0�3	X-@D�-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo�o�o�2_�o�o�o �o0BTf$�<�o������ �� �2�D�V�h�$�������@����$�P �������(�:�L� ^�p���������ʟܟ �Ϗ$�6�H�Z�l� ~�������Ưد��� � �2���h�z��� ����¿Կ���
��@.�@�R�d�vψ�W��=������nCA� �������(ך͚�B�k�Vߏ�B�%@�׮� �߶�������
�,�Р0O�_��DPO�@1��_,z�T`"B�^�}4�� @D7�  ��?����? ���2>���	����;�	l��	 �� X?�X����������, �,X � ����H��H�f�fH�PuH���H�WH-���u�s8��j�|���BO�  B�0����������4  ¾��¾  ��0��������������]�F���A������:@��`U����ix�h�0~&@�  �� �� M'0Т����~�	'� � ��I� � � ��z=��q��@*@0+~1T�;~2��iw� N�0�  �'� �� C��B��0e0�1B���1��x�}�,@�B�L�O���J�dPH{�B� Z&�0f%�:� A�%NADz {ߥ/�/�/�/�/��� #5!/5  '!ȧ :��&A��,>N@�?�ff9�`?<r?? ���?�<�!8N@�?�:��R�4�'(N@EPH/9O��
�
�t�3T1�;���;aʤ;��D�;��;�	�<$DB�DO�1A��j��hy?A ?fff�A�?&�@�$A��E@�,�Ej&" �A���)��_��1_�G ��?f_Q_�_u_�_�_ �_�_�_o�_,o>oo boMo�o�O_!_o�o�{hE�`	��D�:�`�o#E�r�o /zoS>wb�� �����z�#�� H��oi��o�����Ə0؏ꏉK� �?��[!O(��K�6�o�Z���A�A�Ap���  
�ş!���쟃�}E����4��X�C�U����AÁl�D��D��` Cai�V����c�ϠΡ֡@I���COLCC���Ck�B��1B-v�=����n���)���1�W
��u /�R�@���
�7
=AX���Blz��X���2������i�c�ö�=BU7(�¥ ���LJ��LI�JJOޔ�LUW�H�� �I%K�AA��M�DLs�L�]��HP� H��R�������8�LiPJ�
`�H㞀H���A%S���@�+�d� Oψ�sυϾϩ����� ���*��N�`�K߄� oߨߓ��߷������� &��J�5�n�Y��}� ������������4� �X�C�U���y����� ��������0T ?xc��������>)Gj8O%k.D��s�5Ā�R��C�B߾��/��s_�//C9/�:/��/�(r!�`��(/AB���%r%��1V�`�/�-�3Z��b�/�/�"��v�??��v3��g�.?@<!�;�%D93ҵ�Z= Z9�?�?�?�?�?�<�%PzBPN�0�=O@�/IOsO^O�O�L��O�O�O�O;\��O�O�8אt_�Oa_L_�_ p_�_PO"��_�_ o�[�-ooFo4oVkO��Voho  �e 3��oDo�o�o�o��o z  2 �E����7FvD����B����ÐCGpD� A�@ß����Eј F����s�> G� �GED Gt$ ?F� E��/�+[��_�/�A�S�<e��?�ff~��U���T��r���
 l� Ϗ����)�;�M� _�q���������`�	�����+0����$PARAM_M�ENU ?Z5��  �DEFPUL�SE�[	WAI�TTMOUT��RCV0� S�HELL_WRK�.$CUR_ST�YL�\�OP9Trqr�PTB�����CW�R_DECSN(�E�\ү���� �,�>�g�b�t�����િ��ο���SSR�EL_ID  �V5.A��USE_PROG %�q%�X��CCR4���.A	�k�_HOSoT !�!p���e�T%@w��ÐϢ�����d�_TIM�E2�ƀ��GD�EBUG���G�INP_FLMS�K.�]�T�n�_�P+GA�� M�����CHk�\�TYPE
��
���"�K� F�X�j������� ������#��0�B�k� f�x������������� ��C>Pb������_�WOR�D ?	�
 �	k�H!2�F#{AL4�	JO���TE��F#C�OLD%�Z��TR�ACECTL 1��Z5�	 �@C D�� }-@ l m��� � �` � ��  ��� � �⧁,B�~DT �Q�Z5��D � q 9P�	 9$:$;�$<$=$>$? $<p"rp"��"�� "�"�"F$J�*"H$I$J$�Ј"R"M$Ϡ"O�$%@"Q$��"S�$4�"U$V$W�$X$Y$Z$[�$\$]$^$_�$`$a$b$c�$d$e$��"g�$h$i$j$k�$l$m$n$o�$p$q$r$s�$=P"u$w$��$�"#� @DDcpBU!D"D#D$DU%D&D'D(DU)D*D+D,DT%`B.D/D0DU1D2D3D4" ��B��A���B��A@��A��A��A�DE	�D
�D��A�D�D�D�D��BU�D�D�D�D��D�D�D$C�+D3D;DCD�[DcDkDsD�{D�D�D�F5J�D6�D7�D##$U+$3$;$C$UK$S$[$�$U�$�Tdd�$&�C�D��D�D�DT�TTT#T�+T3T;TCT�KTST[TcTjkTsT{T op�"$$�S �$$��"�S�#D+D3D;D�CDKDSD[D�cDkDsD{D��D�D�D�D��D�D�D�D��D�D�D�T2dc!t�#FUTTTTU;DCDKDSDU[DcDkDsD]{D �a��A�0�AM�"M�4"M��<"M�D"M�L#�D��D�D�d�D
�dTSM�T"M�\"t�CU��BU��B U��bU��BU��bU�RU�@�SU�$RU�,R U�4RU�<RU�DRU�LRTU�TS�D�D�D��d�D^�p�Ds�Kt�T[tct*kt�T#D+Dƌ U�\S֟���l�~��� ����^�dRU�lRU�tR U�4sv���������Я ����<rM�d"M�l"r�C��B��B� �b��B�b�@�t" M�|#6�H�Z���0�B�T�f��$6�H�Z� l�~��������ό"M�`�"M��"M��"v�C ���B���B�Ьb���B �мb��R��R�И� ��$R��,R��4R��<R ��DR��LR��r��\R ��dR��Lr�ЄR��\r �Є"�Ќ"�Д"���" M��"M��"M��"M��"`M��"M��"!v��U������#So�C���B���B����B��B��B��C��D�D�D�d��D�dTT
T#T3S��B�� �B���B���B���R�� b��b��"��"�� "��$#������l�~� �Ϣϴ�΄��,#���� ����0�B�T�*4" ��<#��*�<���D" ��L"��T"��\"��d" ��貹�(¹�|"��@����"o�3��2��x}y����+ z}{Q����� @$��<B��DBt�d a `��da p��da �� �da @��da ���da  ���da ��ta ra  \Ra �Jta �Ra \r a dra lra �Ra $B a ,Ba 4Ba <Ba \% LBa TBa \Ba dBa  lBa tBa |Ba lLB ��TB��\C�(�dB��lC�D�D��D�d�D�d�TTT#T C�tC����(�:��rT���������cI�g���@���@�b�@�bn���@���@ �b�@�E�b�@�b�@�b��@���@�b�@�bf
 ��EP��EP�bEP�bEP �bEP@U�b�@xU0U�� �@���@�b�@�c�D�P �c�D�P�c6T�P�c~T �P�c�T�P�c�T�P�U��c�dtt ��@�cV��`�cf��` �cv��`�c���`�c�� u`�c��u`�c��u`�cƓu`sn��@�b�@ r�_�o�YU��O�O�O __/_A_S_e__�o�rВp0e�pذ q0��rز�x(��u�u ����(�5�+� �M�!�z��p "��r"p$"��1 �r$ �r,"�4"��� �r �<"p42p�p � �r� �r�5�r�  �rX�8��p�2U�K� p�2�D��������r�� �r��p��ݓr���r �������p��pL� x �2�vuo�D}� ��}�B}�B}�B}��B}�$B}�,��x�j{ݯ��T�Au������U��������+��i�{����� ��ÿտ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻����� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ������������ 1CUgy��� ����	-? �~te���tm���t m��vTm�3
�#m �Rm�Qh����� / /2/D/V/h/z/�/ �/�/�/�/�/�/
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O �O�O__&_8_J_\_ n_�_�_�_�_�_�_�_ �_o"o4oFoXojo|o �o�o�o�o�o�o�o�0BTfxNow A� B�tUC�tD�tE�tF�tUG�tH�tI�tJ�tUK�tL�tM�tN�tUO�taq�goUw��U����)��q�t�tТ��p�t�t�t*�t�t�t�t���p ��p(��p0��p" �t���rH��pP��pȒ �p���pؒ�p)�t�*�r;�t<�t@�t� ������"�4� F�X�j�|�������ď ֏�����0�B�T��f�x���������^gW Za��g��������ÿտ������������ ,���4���<���D�����L���T���\���Td���������@l���t���|��������������� ���������������� ��������������p ј4�F�X�j�|����� ��į֯���Y���� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?O�yO 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q���$PGTRAC�ELEl�,����_����i��_UP ��������������i�_CFG �똥���� �������گ�ȡ�����DEFSPD� 츬�����i�H_CONF�IG ��V� ��dW��x� �Z�PŤȡv�����i�IN��T�RL ︭ء8l����PE<��F�����ѤV��L�ID���	�G�RP 1�F� �� B�f�f���B7�\)G� H,/�G���Af�gD	�����[��ȡ^�n�ڴ� 	� ��y��ǈ� ���*7�z?����B� ���ϵ́������:����"?�EB=�C�|�|��x� <,1�� ���ߏ������&�� ��5�n�1�~���I��z����i�
 B�^  ��G@�N����;mI���I��p�� ��&��J�5�Z���k������M��<=���������A�L!A
V7.�10betaZ��Y�@'|�{?�^�RBf�x C�+  �u�D� ��0M���@ �[�@ B�  G�B)H5���W� L�P�ѣA�;�^f�A͙����!�@�ff@�33??ٙ�@�Yh�?M�@���s?�����OC��O���?��Ѣ A4�06֫�����-��*SY�STEM* @V8�.3382 H$5�/9/2018 �Ae!@6'����SV_T  �P $CUR__SCRNi�|"�GRO���!PS_SAVE_DOt��z �%Ei�$NO�_RECOVER~�"RESULT�!�   
$P�AYLOADi�V�%_X�*Y�*Z�*�I�+I�+I3AR�M�!1492�"DO��A� �"MOV_'POS@0� 	a5M0�l2SPEED_H�IGHi�4LOW�2ACp��7�3�5�S3e1�!��$k!M��s! � $�MAX_PYLD�Y�70XISINE�RTIA  �n0� �5�"�7L�0�n0�1MOMENT4�4�1_�0SC@z ��1W� 9B?BIN�!A ?BMN�ED\FCLVHPLD�_MODE;BDU_MMY11Y��D�2�Ak M�!�2 � $�1_EN�B�"W�@�A� A�NGL�A� �AAAd�#�AB�A�DCC�G=D�$LST_�@ZB�
$COMP_S5WY��2XY�0�C��1Z/Uk P�4 1�n0P%B�&�/p�/??%?$I=�DIS�!`0k � �S_Gs! | QcZ� #C4�[5�[6�U�4�V�4f�4cqEP�#�1  ��U�r"v���Tv���PMON_QU�Es!��$QCsOU]Q�0QTH� �HO�2�`H8!� I�S�cUE�`�"��PO��s!� $�P�@BUP�0�!R�UN_TOC�^�`DATAs!u���fC'A�0}!IN�DEX$RPROG�RAQ@�0�02?@N�E_NO4t�eITyP4s�`INFOs!�	 �`{]q�2�s�Zq`r
 (^@�SLEQ_NUM�ts`pYP�A�r vH��`SCHK��s � 4�`ENAB|�B�`PTION�c� ERVE?0�y�A܃`�sGCF�q �@�`Jf@�1�b�/$CAR���w��2OS_EDITNs! �� 0PKe1��s$HIDE_r%@Ur�l�AUT�!o�COPYe1�`��,�A� MV�N������psPRUT�B z��N�OUCH�A���AP_PRC{RE�1� l�v`0ME6@IZ�s��`_RSET_D�I)�Ap&QIN_FRO�sN�D.p)��fDSP_Ce@�Br�TCH���A: ��(A�� HSTS�`_�SN�1�!WRN_ALM_�"��G�aF� ����2�IS�q
�@Nz�B�6�����|G��pRGADJs!� h�PX_�0I�q$.P+�<P+�W
)�P)�R)��3�$R�NEXT_CYC���1RGNS�u��0בGO_�#$�NYQQ�EQkRW`O��v��%��!LAރ���)�3SO��u�AT�E�c� IFY%vN�AM�@%��_G>ރSTATU�Pރ~�gMAILTI�̋1E�EV\R�0LAcSTE��1��EL"���p ��ȐEASI�q�2�0��s��q(�!���rOT`A�p�2��1���1�a� ICڲAIB�aQ0E-p�0Vg��BAS�!�ð��UPD_�`� Y$
�&�RM��RԳ0�1�PB�'SSP�c`��&����KS�P	~�� 2 M� Uo0�0��0�e@@� A0���dUŢA��'DOUs��I�k��PR�0�p�rGR�ID;q�cBARS �vۀ�saa��O&@s!W �a_�!W��=���O-P�t �s ?@PPORs�f��C��SRV�)l��~�DI� T_�@P�вԣ@��3��4��U5��6��7��8�џl�PF&�q��`$VALU�Î%���0�1F�u| �u�!*qP�1��(�pAN�#D��,�R\��q�1TOT�AL_I�ذ��PW�Iѷ�REGEN����McX3��c�u�Ql�`TR�*���C_S������sV)�>�:��r�EL�	Хap�2�b��~�V_H&��DA�S9�|�S_Yh�!'R%�S�@AR�P�2 �IG_L3��3UP~�\�_�`��1��ENHA�NC�a T �-��sx񑐝�a��u@F�c]�_OVR�cP}`	ТP��f���rߘv��1��OPSLG3��p���"Υ� �D��J�S,&B]�DE��U�!�f�b`� ���q� �!-�܅Jb�"œI'L_MܤV��p�PTQ�(p@q-�C�UfBV2C@P_h� JMaV1`�V1n2}2n3*}3n4}4n}!���l2}!�@�(Am2IN)VIB�@:' Tx1.$2*(26(3*(36(4*(46( �����S�"�0T ?$MC_F�`� ~0L�!�!�����M68���"�� h�PsR�
@KE	�_HNADD�!!�$$���)CXQ�4=��"� 3Oa�$���!p�03��3REM%2�4I�H�K4a1f8U��e4HPWD � �#SBMS�KU�COLLAB��De�� �� �xpI؝�Q�BNOgQFC�AL�B�%KT ,�^@FL�@�$SSYN� LMPC�����UP_DLYz�A�bDELA=@�J�)�Y� AD�Q�Q�QSKIP�E� �v��`O�@NT!��g@P_�`r�G pR=��G>��I���I �ЪJ�ЪJ�ЪJ�ЪJ��J�J9��JS2Rs��P �sX�T��LQQqq�LQ� B�LQ;q AH�RD�Cw��2! � DÀ�R�`� "!RN�p�Z�b�R��RGE'�8ó�S��FLG�a�0�� SW�y��SPC�Ps{�UM_LP�2�TH2��`?P 1  ��	�v�p11la" l� `1�0�s�3ATC0 ��� 瀤vfb�p$t]a�p��\b�c"!HOMQE�b�/d27b#=o�Ooaoso�o�o��0c37b$�o�o�o�oW l/d47b%7`I[m� }P
1b57b&����(���g67b'1�C��U�g�y���&w77b(�����ҏ�����w87b)+�=�O�a�s���� �S�0�q*  �̱0c���PcAa2E��+J �P?���&=�IO�]�I�i�� :�R�`WE!�, '�
@jQ 9/`�� -E��$DSB� �g����8@C`i�?��RSw232C�. ��P�0� ICEU��E&`q�PARsIT~��OPB�0�p�FLOW��TR`���r1��q�CU�=M��UXTA�0q�> ERFAC�R0�UD� �RS;CH�/ t� � 6\�EC�S$^�]�OM��A�Ph�IH�##���A	��T�������@̸��� E�FA6�"�1RSM�Fg���CK 0� L��З���M��Ű�E{�x�NSE_*�!D��Y�A�B��A.`��CT�RL_ 1u@ȧ���A k�FF0�����|�PX<�'��_���GPMV�$?SEGFRAp0"
�Q��Mh����U � �20 ��P(���?PO��T����C�) J�5 J���DIO�2 E@~�a�A�֕��V�3D ��DS�3��˰v$�_DRX@����A��Զ�C |¤�ùO��x�D�02$��AL ����INF��_HAP���\��h�Y�AJ ����oՅ����+�Ε"ITR�̒Z_�OFF��	PAU�S_� 3O�r��$7MNT�CMe3��T fUv�6�c�4� 3���4�� ��� �Q������CHK� ?���/�`� ���QCOU�REG,�eALAM�P�D���q�SPG�ն���B� F����2ŢV�`��[�5�˱W�MO�PsOU^Sm�STE^S����S�~�DI_���J���m�OPT��U�PO��
�	c�����6�����0EC�5 8IP!�Q$�(�DZ�OG72�t`@CDI��� 6� D $U��M3SG;�SBEVB�Nچ@�ED@��(pE S{HA?S7 <IQ�*�<���)Q��)Px�P<d�~�8� �1�����A����PEX`�IOE1Ѱ1��s������2l��WR�0Ο��D�Q��P�OFRIEfJ�U��yME��TOOL��MYH� I�LEN�GTH_VT8�F#IR`�#�P��Ѡ�*)U��V_-p�@�(�RGIWAITI�B#'X�A2)u&G2uG1~�oď"�'P���cO_ �����0!Y@�P�4F�{�TC�01"�!�&�M�G�0m�~�9 @� �P����*�j�8�j��A$��0���6:X ��M�C �"gP��P/��a4GcW���74�Һ4D[@LOK �4@HC�@��1�4�A��4 29���7`R�1�?�2�2K3�3�IeA�,I@�A�hM3hY3V�J1"Vv%V�@1!l1�"�;�Pk��3�@�&C��K� Zp��PE|R0#���$4XPRfP6VL5Y3S�@ơH�8�4F��< 0��`6@:� �D@;���G಑O  
�5S��/= ��AR������ ��N��AX%��0A� L!\��RgTHI�!�LIշ>~�FEREN�Q�U#IFG ��QI�6c��PG1QXUd� \iiAf!�tf_J���ePM�P	�RTD�> �젪�$����B�1
`C+��`� U�!���D�`�w�INWo 5�$�TBC_P CMrw�D�aʶLDR���S��&q[�Q���S�WITʒ8���ATEA~�?<�\p�� �a$VALUqq��Xv��e�@��\q  2�? �SC��A�	� �$ITP�_)$���sTO�T�T�su��vJOG3LIL���_P�0B�1O�Q*��AX% U�K�MIR�q�� �M|20�AP��81E8�ʶ%SYS&� ;PGe�BRK�"˶�NC�PI��   ��Sӗ��r�a��s)�GBSO�s?�NÅ�6�P��V�� ģ�FSPD_OVR4 �P�LD���COR�Ɛ���Fal��pOV�uSFB��PE��F^�����#�v��V�LCHDLAY	�	����0�pW`��䷒�pROA�ρ�p��  @PY�I �ER��s���yp��WD��"�ρYI��b���!F��K��ap�B*��B�d���@cTV�������s>�9��Dl�AMh��`����ג��_Mn�N�����T$CA�p��[cT$HBK��ʶ���5�T��I�PPA�-��=�%���%�~�DVC_DB��@n���o�����1��$ף��3��ݐA��f�0Qo���U�*p�� AB��:���J�x��q��p_AUX��?SUBCPUf���S�S����M3AǜY3��FLA|a�QHW_C@�p�3s��3�A�!�P�$UNI�T������ATT�RI������CYC̑���CAӲ:�FLTR_2_FINd�TART�`� شB̂�LP��CH/_SCTG�Fe���cF_��&ү�FS���Ҙ�CH���g�b�r�RSD��*p�g�v%�_T��PRO��.�pEMP�P�p��9TTүA TҸA��Ւ G��RAIL�AC|�@�M�pLO ��#ۄ}�o޵}޴fףPRp�y� �PzE�Cb� 	֓�FUNC�R/RRI�N0t��e�qRAv�� ����2���Ύ�WARmc�BL{���A������DA��������L�D��1!��q��p!�TI|A�+�P;$g0RIAJp�AF2�P� n�ϐ`r�+@�2h�OI���1�DF_ ғPD�R�L<�A��HRDY�O8 q4 �|���MULSE ���A��A��J	�J�$�9�4�FAN� MsLV��@WRNG�� D� �Ay��2$� DOW��[`Qa}�
�@ STO�rx�_���AUx�(px�� O_SBRd���p��
��d�m��MPINF�P����gREG<f�DGP���#V��Y!�>��87����qB �@��$�$Z�Q���r�q�pC� ��]�EGI��s�AR�p��2!����j�AXE�wROB �z�`�v�a��_���CSY�����	&S'�WRI���s�ST�R�u۠���E�Hvp�Y1���BS ��Z&jQ�àOTOrvp�ARY�s`�"�ô�q�FIs��$�`K���Q�!%�A_P#��qQ��"XYZe�*5N�&OFF됰"�"J�(� B�pZ�640����^�73FICP7ЯQ��Z��t_J0�qtr��e$� i$Zs+6�US��B�1d��2C��Y�DU�º�7"�TURB XH��5�!�X" �7FL�@���@�%�V*8��� 1BJvpK�MĢ9"�pA�I�A��ORQ���q��X'3�>�p�i`���J��E���q=�DOVE�A�RM�ha\ �Eb�Eh�Ft �Hq �G��Dze_��s��Q �A'�;P��ha�E�A W`�Ub�U S�qER�q
��	&�E��\p2��T	AqQ��S5��ҝ' ��� �AX��tr � -q�ѳ!e��)i)i � (j0(j�0(j�0(jP@(jv@(j1�(f�� %i��5i��Ei��Ui�� ei��ui���i��i��x�i�a�iDEBUk�$f�r��fq ��"CAB ���&��CV�j� 
�r���Q�u [��w�!�w�!�w1�w �1�w�1�wPA�wvAx�p�0r�YR73LABM2q�Eg�t�GRO��4�2kܠB_�ѪV ?$�G0� ^����E�����ANDd@&��T ݱ�%�Q�ׇ ܡ��!�������� NT�R !��SERVE��wD $40��A6��!7�PO�o0�9�� >�m(�q�v�E  $[�T�RQB
Z��d�F�h�r�2Ey�P���_ G lP�����ERRs2p�I�V8M0XS̑TOQWTTPAL�'d/"ߖ��G9�%�! � lZ�� c�GH ,5�}���F[Q�RA!� 2G �d>�%��p� IW$�@�Ң�b�,�Z�OC��d�J�  ��COU�NTS! ����S��rK� �mM+�>�hPEL3AY׭�VAT*�G ���J���M�	٣#GCSFs0P �K�À0�b.�h.�׳0�V�+�.Q �FX��m�YZx�Zx�NU��V��Wx�HP#�
�aƲ ��ӴbݷhݷV�ݷpa�ݷtZQSFIxp6	�IGQ�DO��#���%�܄#�x��Q��2���L � �?�bN1J#��4SF"�Q���2�FZN_CF5Gc�Mt�$?�T�L�q	aZs��R�� U{�����N ��pMh��Qi00SS�Ah��FA_�bUm��X�:�����R��:�$NE�P�h����DS_PT oO ��pSPyІj�DU� ��m��D%I�40��Ih��&��SE���W�Л���$DR�Ab�0B���V�mHEL�L��P 5�0B_BASƓRSSR>���S�:�7�1�7�2Z�3�Z�4Z�5Z�6Z�7rZ�8�*�ROOš�%�!� NLb�3AuBF�6�ACK�v{INl�T_CH�1�  � ������_PU��1lS�OUH�PN��AA� �	���gT�PFWD_KAR�ё�p��REE���P:� N�QUEA��P(�@�0�C�IC �s��� H��#�!SE�M�q��c!���S�TY��SO(ċpDI�� S���g����9MT���NRQ6� ����C$KEYSWITCHH����HE�0BEATmM��PE�LEВ(��z��U\�F��]��SDO_HOM�+�O<Q��EF�@PAR<1b�@ �C� �O��E!�OV_Mx�2o08�IOCM�4d��c!���HKvGQ D�!C���U��£�M�w��@�3FO�RCG�WAR�� �  ���.�R �@ptl3��UF#PA�R�����3�4��� �q�Om�L�S*�B�UNLO4#��ED2��@?�SLCL>Ac��Tl �AN'CELH�*&I4%���DRY3&J$A*WETQ*n A%����3%�$<A%�ZON13%�%��,2�,2�,3�,3��,4�,4�,5�,5�A%�k�3%G4A%PU1R7�^9A%SE'���x;w6�Q�B�9w6��P1�6�4�7Y��B�7�3A%RS�@�3%�5:A%U8�DEF�&E L�&=EL�&]EL6�}EL.6�EL6%L6�L7%L7L8%L8
L9%L9L�P7[w6�E�&]SUZ�&ySUZ �&�SUZ6�SUZ.6�S UZ�F�SUZ�FcUZV !cUZ$V=cUZDVYcA"?GI_BCK\�Ѐnlme��zh�eme��E@zh�e�f^W�fA#O!��7�g�fT��fs	xe8-w	xSVhKy�eB��H_RG�lx�e?CLR_XF��|�vYC�^�y�ez�|�eЯpLv�u�w �)���$-���$M���4m��.4���eMAJ��p$�����s����s��г��H1AU����? �? ��BY�vK��T_N0C��m��eNO�!�����ePOWm��5��<�ek�T_RDP$ɗ �e2���e��eK	� �6�MK	�V�mK	�v� �K	����K	��D��� �Dɧ�T��$T	���vM[O_{��K�C�4 PLr�k��^X ����6��Y��V��Y�� v��Y�����Y�����Y ��Ҧi���/i����Ki���vgimpCKP8�&�ț�EQ_H���Û�FAUQ��ś�@���'�ț�Z�qD����DA��9՛��� ��Y�Q��h��-!�x`" U 9B��`x`GROU�LAST_BIT \
�`ERF�!E��Ƨ$_T6�Yb�INF H���@I��B��O��p��"V���&�S�sM��(�E_/WIDTd���SIZ��ːl����q�����TP�p0  c�i FIG��(����opL���ӻ`P������3��4
��TO��  	�e2���AIR��F�h�Q��e24"EF�� P���3�TO�G��k�CC���3G���SPX��o�(�m���l���l�5i�6*i�7i�8i�9i��� ���������������� ������������������\`��N(Z�� Z��Z��Z��Z��Z��Z���!��>!!V  d��F  ����I�SCFG!!W �� $!D��H�AN����J_CT�RN�$IS����T��IE(PD)S�A)��VO_TY/PE � 	e��Bp'6�тG��W��MB_HD}D�� X � �BLOB   � �SNn�AS��Y 0 $A�DDRES`�$�M�$VAR_N�A�%$M��P�LYW���A, �Z � $T�IME��$�_I>�	$��7"��CI2�Q#FRIF<7"�`SIONa\��U��$6�INFO�7"G0BUS_AD�RN&�#�)P��U�4�SPl�TSK~��[ D x |�a$WLDr��$XTRA_S�H��u�$��_M�SK�CL� ��\��S@� \ x ��NGLEST�E��$DUMM}Y��$SGL+1+TA0�&x D3�<1,0STMT<l\4PSEGl10'BWD+6� We5SЯ�SVC��G��] ��$PC�p���0��	$FB�r�8ScPC[�7� VD�0�R��^� �]$>�A00pt��21�92�93�94��95�96�97�98��99�9A�9� FC��9D�9o FF�81��91	I1I1#I1�0I1=I1JI1WI1�dI1qI1~I1�I1��I1�I1�I1�I2��92	I2I2#I2�0I2=I2JI2WI2�dI2qI2~I2�I2��I2�I2�I2�I3��93	I3I3#I3�0I3=I3JI3WI3�dI3qI3~I3�I3��I3�I3�I3�I4��94	I4I4#I4�0I4=I4JI4WI4�dI4qI4~I4�I4��I4�I4�I4�I5��95	I5I5#I5�0I5=I5JI5WI5�dI5qI5~I5�I5��I5�I5�I5�I6��96	I6I6#I6�0I6=I6JI6WI6�dI6qI6~I6�I6��I6�I6�I6�I7��97	I7I7#I7�0I7=I7JI7WI7�dI7qI7~I7�I7��I7�I7�I7�D 	X�0PR��G� �_�|��� 
H�0�"�!`� $TORG�0�D�� 䩠��E=�Q_C�URRE�2��AX�'���� YSLO~�a � ���"��y(�� �0L�$��2VALU�OP҈�$Ρ7�F�ID�_L�#_�H�^�INFI� n䋳$�$@! � �S�AV�!b h 9$����LCK~#ò|F1̸D_CPUܹ�M�ܹ�Z�������Y�+0,1 R c � PW	�`=�	L���R��_S�L�RUN_FLGe�.i�L�WU�mĊ�.Ċ�L�H,��L�U��TBC]�k� dX -$���LEN��������EgL_ROЌ!$W_ܡZ�1��w�2��MOԱ1 ��E ERTIAդ��8٩����M�DE]�6�LA7CEMӧCC+ӵ�V��MA�\֖�l׎��TCV�ܾ�l�TRQ�������2[�sH�l�sJZ�4M'�"cJF��0[�H�l���2'��0� a�Z�6��JKt�VKV��xc��p$JJ0�䶊�JJ��JJ��A T������}����N1����ۚ���yL6���H����e `��GRO�UE�G1�"�1NFL�I�"J�REQUI9Rà�"EBUM#��n(�$T��2d�����l�����3f ?\ $EN�/APPRx�C!�п
$OPEN��CLOSE���� c ���[�
��!&g �MC������_MG��) C�0��3�(�� 4BRK2	N�OL�4�"MO_CLI�!xb#J� tP��xВ�xК�x���x���x�6�91��0 �Ţ�h� u����#��PATH2(2���.# ��g�О1S�CA��x��(INF��UC<Џ!�C�0UM�Y�A#�c��E������D P�AYLOApJ2=L�R_AN����L>����
!3R?_F2LSH�"4$LO��8'�F'�ACRL_̱�x ȁ���H8���$yH3�"FLEX���+�J��i :���ư��'�$�ϔ�0������F1�!<5 P7&�8�J�\�n߀߀2E�ߜ߮��������� ��WHtD�3�t�d0@�H;�M�_��!f�T�GUAX�^Ar��4�8}� %U�8��������债���������*�J>0�j � <�N�`�r�ATi6t�&�CEL�0��;c{�Jb�i��JE_ CTR��d1TN��7fl�H�AND_VBB��!D�k $�@Fa23��QP3�SW%��l� $$M   	��O�h^�l@�e�vAf��#e�D3y,A=(�O
A]AAl>p>��O
D]�DlPLGT��yS�TQ�q^	�qNoDYk���3tFu �� .'�!.'I!�t�D0�@sP�����������"m �`�$��ن���ASYM\@�u�\l@wI!|_ ��m(���+��h�����J�� *pʓ��*)v4_VI�c�����V_UN!I>#,�NS6!Ju�E� s�E�I,I�`%V�z�i-�&�|)� �/�/ͥS��$�#UŁCPPI>?� n  	����@Pj� TCDEwLAYOQ  ����SPEE�  o# X����@N��RP+���� M�����E�t�1(�M��$PR���V�q`YPE����_�0�p |��"��S�Ep��S"��3fWoARNI\�EN�`� OTF0�ֶl�_�T�U�MA���C��f+�CP_HIS�T_BU_ q� ,�@P`2gPR�z��U� ��SPD���r ��P��`E�ARTBE7�SE�T�P��U�Pp AR9G�l�FLG�%�ò3S]��TR����Ǣ���I!�#�ǽ�R�E���NR$�`�OU�T�!s p���T�E+Љ�r�B�ID�P_$ʠUn3+d؈�K�Ju�׳�S���H�����t�b���In��$DO�� +�Ж�u ^PMrI0�A�|����U����0G`���1��vo � �aME�1�g�Rc�U�T��P"V�D��!������J�e�Y�T��"� �$DUMMY1�VQ$PS_g0RMF)0  9�� �FLA2�Iպ�X�GLB_T�`׵�������[��0ha��w5��k�ST�1��S�BR��M21_V�[BT$SV_ERb O���3�CL��"�A�0C���D��wx �(�TPS�0��1xa*�ADN��$FORCy�BA�CK_FIp��B�GLVkc��1���v�SIZ�������a�CANAGE�_ME�$RE�CURSW�$AH Wa ���NQ܏���PGL�EW��!y 47�Z�$�$ZORWQ�4 2�cA����[�3]U7z �@Nk ޣ�$GIx`}}$7 yl1j �!{ L7����)}����E�N}��0�Nn3F�	�0TAN�Cn2��Jy�R3q �|��$JOINYT�@  1M���!}��E��1`�Sb�`�!~׼ e0U�1?�@�LO��O
곫��GL��Tl�_XM� DEMP[Bn�x���p$US:�8 002z@�j�{К�`u�y@�CE8�P�� $K��
@�M��_�: $VE1C� &IU����CHE��TOOL�03C#V/4RE% I�S33a$6�Q��CiH��\`}P!ONV�&��29��Y I9� �@$RAIL_B�OXE�@�RO�BO�?�@�HO�Wϱ�$���!ROLM���%�Q�$�"�Q �X0�`O_F�P!G T}!���u ��u���SL9O0 �)�	���y��Baapu�IP�N�@Y"�"`}!�P�00��OR��u\`O00�PO� �� D ��OBsqEcu�7�1�㱰��2��GaSYS�1AsDR���TCHpG �-�6�	_��>D�QL�uVWV}A��� � r�x7׵2�V_RT���$EDIT�FV/SHWR�Q��@sIS� v�IND/�RFQ�DNQ{�D��hǠ�@���CKE����^��FJMP�0LLֵ� RA�𖴅�0U5�I�SFbC�`�NEL Ga�gTIC)KM#:�M�Q/S{HN��� @�0�1Q��_G���&��S3TY:҉!LO������R}R�P� t �
?%$cA�=:�SY�!$;�M �4�I���H�P��VS3QU���LOJ���TE��P2���T=S��� � �D3nbD����m�T:!t�OJ�=�����GՉ��w�C��b۲U�TPU2��e_DO��=@XS(KֶA�XI�`	3�UR�U��$T� oP�6>:�FREQ_: B�ETrP~�0 ���PF ��P��DA�����#�#�� tS=R˄�lO`�� n�4�+��r�z ��~!Vb��v/��xAY�	h�ww��|AˀAV}� �u�r��q�D�~��"�D�� �Ce���C�z�������a1S�SC�� � hF@�DS�ԏ���X��AT��q��)�;T��ADDRESM#B��@SHIF���_W2CH@�1I��N��TVZI�ҋ�-ª��H��`
�
���Vh1�aj�� \��8��P}�ma:��C@�pb3r���69���TXSCREE��2����QTIN!AV� ��tq���� T#Q6��� Q��Z��aB�b���@RROR_�E�R�����UE��� �`�p'A�� ARSd�<��׵UNEX9`ֶġ��S_d�~cԡ��~cqCj��A�o 2��UEqs����F�'�w�MTCN_�����"�O���BBL_� W�v�j� ��P��O^��LE@���� �TO_ㄱRIGHΤ�BRDH�6�CKsGRv�̵TEX�`͵ȱWID���@�7Č��M!��U�I��NHz� �� 8 $�T_�AN�+�/�R�@p�#���u �OG�j�xPS�ŰU��y�R~�!LUMy��f0�WERV���P� ��i�&�DpGEKUR�F.p:)�@�LP��,rE6`��)���с�����w ��5*��6��7��8��4b@|c�`� Δ��w!h�S:��USR�7� <�.�U8�b��FOC:!� PRILqm� }a���TRIP�!m��UNDOe��� `�P�����!��X��p` �&ОaG �PT	0��O�&!�OS��6�Rp���I!i�@RY]�H�T���U��i�f��x����U�OFFT�j��0��O��� 1�@�����N@�GUN��%PB_SUB�RO�=�'SRT_�qt�xR��0~cOR� U�RA�U�pV�Tk�&W�VsCCƠS� R1C36MFB1�d�  \��p��Gx �"�1
ci���a���C����D�RIV�fq_VЊP��JP� Dv�MY_UBYu����V��`%��A�Si!�P�_S�0coL�kB�M��$<PDEY��SEXq���ia�P_�MUPX���٠UASQ0�2��&aGܐ�PACINLQ�PRG�`����������RE@�D�I!$�����`���TARG P�8=�r��RM�-0� dq���a�5�	��aRE6�SW� _A�&�I��`O��6�AH���rE|`U�P�!&�YfP��HK�R�xP��'`�q�_��E9A^P 'WOR-���!0=MRCVD��� ���O�PM-�C��	="��5="REFp�_&F&1!���=s ���B*�!S*�!d+�%F&�_RC+�(+�0ScЫ"_aha<�=A�� ��R���p�0��'@ROU�Wx0�V�� �O��2�K��А�`LP�����8RK�`S�ULA����CO���@�� �0�C]� �3�A�6Z��6���3�0LY
Ei
EZ�G������T�t �+�EqҀ �CACHcLO�!]DsA� xI��ZcC_L�IMIA�FR�HT8�p�F';$HO-��R=a@COMM�����O���GP8���VWV�P2�QQ_SZ3d�3&U6C&U12[�`#X� !X�@!XWA�E�MPeZFAI�@G��r@AD�Y�I�MRES4�R_�fG�PƠ� �p�ASY�NBUF�VRTaD�U�T�Q߳OLI�SD_��eW��P��'ETU��@Q��U�ECCU%VEM�\EWb�GVIRC�QeVT�`�e�b�V��Sr�Q_DELA@*Α�f`��A������CKLAS#�	$AA�pG�Q�ҏA�S�PnFNt�LE�XE���M����,��FLɰI� �SFI`Hw�0Gx��C (!�aRpE���-z-4zԂ�]���7ORD��� z��Ш��Z2�����T���[�EO���s�V=��թ`�0F��@�UR��_R�P�B���ST� *o���@�����x���T�p��SCO>���C?�� �� � �� ⺆ �Ǉ �Ո�������K�Z� �EڰAiM����;SM�����҄�$ADJ��p��xQC��8���w*�LIN��������� x�MGSPD=���R ��`"堩�LNTʣ��M�pA��g�Հ_ACCg����'2^$$ZABCB�����Z��s~ 
51ZIP��ծ��DBGLV� SLN�~ ��H�Z�MPCFB��  ��Ы�ۤ��1LN�K$�
X�M�C��� ����A�e�0MC�M� C SCART�_���P7�{P$J��DQ#�4��-��9���UXWM�¥UXE�g�b�(�_�>���p���p���� ��Z��g� ��N� ���uYǐD� �&�:I���IGH��x�?(�0ǖ}!  |��>4� � �t,j!x�$B�0K�0cK_��3��RVi`qF��~"�OVC�����4�p$tѐ�
��"I��UD��TRWACE�`V��Ⱦ��SPHER
  �� ,�0���"� ��$PLID_K�NO�  ��-���-��SV  ���J�{7��-� 
 -�m�ߑ���  	e��ߵ���B��d_��
�=�M�ac 1X�L��@�B�p���-�������^���@�qd �H-�@�-� p����� ��Ѯ;3 1(�T-�Aǐ  9�9�-�C-�d�B�����l�xњ��1 1J��U����4T�ool Chan�ge-�A�p�V����b��B���G��G�"ߟG�"1��� L `�& Pa�rt-�B�  ?���@ p�ffG��A IY�Ix_�����Only-ԭB��?����.�� HT]�Hty#���274�������\t�T�����#B9X_H�h8G�Z�G���������B�[����q��F��8 H� H{*r��311�������bt�Yk���U�sB4q�H�?�G��G��2*d������s��������erBB��H��G��>Gw�;���336���AL��ܓ��y�A�B�J�l�G�|�V�� ��A��t�����2���B�R���v���39��t��G���l�B�\h�k����h��؁-��2 �q E��A�z���:���Fm�B������u�b���\)��H�RXB��fE����D��7?3 ONLY���R�#(a �r��q^  녢��7\)G� H?,/�G����� y�k/}/�/�/�/�/��/?�/?R?6�P2�J�\�;? �<�?+(?�3y?�?�?�?�?�4�?�?�?O?�5 O1OCOUO?�6rO�O�O�O?�7�O�O�O�O�?�8_*_<_N_?�M'AD �`�U�7OVLD  M��W�^?A��̑ p�_�:o8�SCH�Z �UTg̑bi7�teUPDo/i�o�d?�_C�����PK�Z�'q5��d�CHK�e��5��b�o�k؁ +�=�p�DVw_B�5�_RE�I�M� �r�C��qB��H;���qGi:4o�_�(+�C��S�B��{H�u "�G�����w C���=V�B��9H�{2�b�G�Zn�ޫ C䲏v�Bֿh�I 傁G���x��L�C�-����B��-H�{ ���G��W���C�����B��qIvG�̗���GC����ցB��I {@��G��.��@��C��\�By�
Hܶf"��G�����C��T�6�B��rI� {B�G��� � �_�d��������� ݟП���]�sx0�|��Q�%��r�0?�^� c��s@~������sq@ ��ܯᯗs�@��� � �sP;�Z�_��sjPz�x�����rV 1J�|1�4��T�pXr?THR_IN�!�d5�d�MASS6� Z.�MN�L��MON_QUEUE J�5�cp:�U�4N�`UqN\�{��END�����EXE�ϻ�`BE� �Ϝ�OPTIO��ǈ{��PROGR�AM %�%���ؿCo��TASK�_I�T�OCFG� ��_sߦ�D�ATA!����@��7�� 2 tru �m�,�>�P�`�t�� ��#x� �� u��K������%t���@�������� �0���IWNFO��	�ݘ����}����������� ����1CUg y��������5IK�
�� ���6[`K_����k��&G��25 �P(O�=����w��@�  � ������!_EDIT ����ڿ��WER�FL�� �k3RCR�EP 5 B�����L!' 
��q/��y/h6�RGADJ ����%?���%!��&���0�f�;?�L0&������<���k�%DIAG�/4?�f	��%���2�V��	H�pl�f�"Bp�� ���@� �=�*�0/�2 **�:�2�?�6CM=��`"��R*�4P�� �0�?�0�/O6HC�*w  F�1����bmPn�ʰAC��9O.O|O�KD���L@���TJ�pdF�UUVpO�O�O:L��؆`���,"�f����O�O__Z_@F����`�(^~�dF��pH_r_�_:LS��`B#p �֡sagAʰk���_�_Ri$mo o,o>o�o�oto�o�o �o'�o�o�o� fL^p���� ���k�>�$�6�H� Z�׏��������ƏC� ���� �2�����h� z�������ԟ��� 
���Z�@�R�d�v�� Ư����Я�_�2���*�<�N�˿�� 	 �����μ��ĺ������FLB���,��ĥ����%9_W��t$ \��J�Wl�W�ο��#�����%PREF' �*���!;�RIORITY+���ր"!MPDSP)�/
�UT�֊3�}"!ODUCT�����ϡ&OGe0_TG 7��I��TOENT 1�� (!AF�_INE4������!tc�0�����!ud��!�!�icm��J�XyY�#W�  ����)� �1��������������� ��	�F�-�j�Q����� ����������*|��#��� %HOM�E_IO 1 C�I�ϴ�=���<?Qp;?+z�3�2022/04/�16 10:45�:305-�����E8H9!dA2,�  ���B�!$���N{���A��6��Bo3J�T��U�ENHANCE �)9#0�A�%ɿU��������E�PORT_�NU�P7����"!_CART'! |j6��SKSTA4׻ �LGS���j���0��Un?othing�_/�q/�/r�# TEMPG j�/�5G �_a_seiban���/2�?(??L? 7?p?[?�??�?�?�? �?�?O�?6O!OZOEO jO�O{O�O�O�O�O�O �O ___V_A_z_e_ �_�_�_�_�_�_�_o o@o+odoOo�oso�o�o�o�o�)VERS�I�V�p �disabled��oSAVE �j�	2600H�607�h�oo!`nq�"� 	�xH>�ÿ�{���e� :�L�^�p�~�)��豏P0u_�� 1�j�\p �;����������URGEAB����6�WF<�DO5�[�#�W��]���WR�UP_DELAY� �P�R_HOT %�A�m�ݟn�R_NORM�AL��r�̟!��S�EMI �&�e�'�Q/SKIP܃��x�o���oί��4� |�#��G�Y�k�1��� }���ſ׿鿯���� 1�C�U��eϋ�yϯ� ���ϙ������-�?� Q��u�cߙ߽߫߃߀�������)�;ￕ�?$RBTIF^��RCVTMOU'���Y�DCR�܃!�� ����E��(D?f��E��Ck�sB�m-B�����R�nŀ�}^��J�.� (���᭵���� ;���;aʤ;�D��;��;�	�<$D�� �j�{� {������� ������1CU�gt�RDIO_T?YPE  �[��qEFPOS1 �1"�
 x�Home Positio�&h\̀��X�X"����?�����`�����6{+�<��5,?�5?�  D́�Ref/Po7unc�#2ʇ��	��0>�rU3f�x/���
Z4f��y//&/8/Z5f�h/�/�/(�/�/Z6f��/i?@??(?ZQsk�X?��?|?�?�?Z8f�@�?YO�?OOZ9fA�HO�OlO~O�JV10g��OI_�O�O��I�2 1#�� � ?_�Y� ��_R_h_<o�	3 1$�_�_��_�_to�_�ooS4 1D�:oLo^o�ox%�o�5 1&�o��o�o�o��@S6 1'W�{��3��T��S7 1(�(��"�ȏF��>j�S8 1)���������]�ۏ~���SM�ASK 1*� p� ��ʖ��XNO����u�MOTE�`���_CFG �++�(Uu�PL_�RANG'�c�e�O�WER ,�����SM_DRY_PRG �k%R��Я��TART �-��ުUME_P�RO����:��_E�XEC_ENB � P�k�GSPD��U�]���l�TDB�x���RM����IA_OPTION~����5�INGVE�RSݱ�	�)��	I_AIRPURn� �NϲMT_��T��)�s��OBOT_ISOLC�L�+U{��/NAME��ϵ��_ORD_NUM� ?��I��H607 .�CVL �rodv(�cs �etu �w
PC � pr ����u�PC_T�IME{�g�xu�S7232D�1.����LTEACH PENDAN}��@��H�'��AMaintenaM!/Cons������"��TNo UseH�����!�3�E�pW�i�|�NPO��f���y�CH�_L�/}�I�	����!UD1�:���R��VAI�L���3�SM�FST_CTRL� 21� D%9���� ������K������  Q���/ASew� ��������� ��*N�}� �������&/ �J/=n/]/�/a� �/�/�/�/	??-?/ =/j?9/�?�/�?�?�? �/??OO)O;OMO_O qOG?�?�O}?�O�?�O �O_�?�OI_[_m__ �_�_�_�O�O�_�Oo 	_:o)o^o-_�_�o�o �o�o�o�o�o�_	o6 oZMo~m�qo �����+�=� Mz�I������ �O��'�9�K�]�o� ��W��������Տ� ��*�����Y�k�}��� ����ů��՟�џ&� �J�9�n�=�ׯ���� ��ӿ���	�߯�F� �j�]���}ϲρ�� ������)�;�M�#� ]ϊ�YϮߡ������� ��_�%�7�I�[�m�� ��gߡ��������� �:�	��i�{����� ������������6 )�ZI~M����� �����)V %zm����+ �//'/9/K/]/3 m�/i�/��/�/? �o/5?G?Y?k?}?�? �?w/�/�?�/O�/&O OJO?�?yO�O�O�O �O�O�O�?�?"_�?F_ 9Oj_Y_�_]O�O�_�_ �_�_oo)o�O9_fo 5_�o}_�o�o�o�_;o %7I[mCo }o�yo��o��� �oE�W�i�{����� ������6� %�Z�)�Ï�������� џ���ˏ�2��V� I�z�i���m��ͯ߯ ���'�9��I�v� E���������⿱�K� �#�5�G�Y�k�}�S� ���ω���ѿ���&� ����U�g�yߋߝ߯� �ߗ�������"��F� 5�j�9��ߙ����� ��������B��f� Y��y���}������ %7I�Y�� U���������[ !3EWi{�c �����//6/ �e/w/�/�/�/�/ �/��?�2?%/V? E?z?I/�/�?�?�?�? �?OO�/%?RO!?vO i?�O�O�O�?'O�O�O�_#_5_G_Y_/O�$�RSMFST_S�V 3�����Q�a@�]J*�T�O�_aB&TaD�Y�Q�]�aB<@o�S�RMA�SH_ENB  ��] �RPRG_ALRM  �[�
�O�oaCQfDSBIL=`�UIn�Q4@n �Q�\�i�Y�e
�_�b!u&x�U-qAvo�h�_CHECK �5�ocwMNCON��P?nfsDIAL/M 26�[�@�_p�y��xfsRUNY`�M��uSHARE�D 27�[  ;AaEF�X�j�|���&��TRB��vPAC�E1 28al AO�}}���R,p�qk)�8�?� T{L�T0�����z��� �������ȟ>�`� R�s�6��������U�Q ĭ�������>�`� R�s�6����������� ���Ŀ:�\�N�o� 2τϥόϺ�ܿ� � �$���H�j�l�.߀� ��xߊ�������� � ��D�f�X��|��� ��������
����@� b�T�u�(�������� ��������<�^�P q4�������� &8JL�0 ��z���� "�FhZ/,/~/�/P�/�/�+ǅ2Ў� �//�/</^/m?�?@Q?�?�?�?�?�+3�/ �/?#?5?�?Y?{?�O��OnO�O�O�O�O�+4 
OO.O@ORO _vO�O �_�_�_�_�_�_o�+5'_9_K_]_o_o�_ �_�o�o�o�o0�+6DoVohozo�o: �o�o����8��M��+7as��� W�������4�U�<�j��+8~������� Ət����<���Q��r�Y����+G <N�� ~��
�7 ӯ  ��� �(�:�L�^�p���ۘ�������d���d ����)�;�M�_�q� �ϕϋ����������� ���ϗ�Q�c�u߇� �߫ߡϳ�������� ,��1߷�q���� �������������+�w `� @��d�̿r�N�V���� ;������������( :X@��^h z�����H Zx.`��~� ��/���
��c/��+_MODE  y��y)S =��R/����/�	?.:	)?R?s�CW�ORK_AD�-��W�AR  ����0W?�0_I�NTVAL� Д���*R_OPTIO�N�6 �%PTCF��>�-�>4��(��,C�2V_DAT�A_GRP 2@,�詑DJ�P??nO ;?�O}I</�O�O�O�O _�O+__;_=_O_�_ s_�_�_�_�_�_�_o 'ooKo9ooo]o�o�o �o�o�o�o�o�o5 #YGi�}�� �������U� C�y�g���������я ����	�?�-�c�Q� s�u��������ϟ� �)��9�_�M�������$SAF_DO_PULSt0��+��C����CAN_T�IM�!Z��5��R� A������@�@
��	%2�!��!��K� �O5�G�Y�k�}��� ���ſ׿�����(�+�226�d����A�M��K��!�!g�O�/�χϦA�������P��2"�/_  B�CT�0����"�4�A�T D��A�j�|ߎߠ߲� ����������0�B�T�f�x����%w���
�������z�PA;�o�D��$p��
�u��Dk'4��+�X �2�!�� ��	���x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/�A���q/ �/�/�/�/�/�/�/? P/$�-???Q?c?u?�?��?�?�?�?�1?�B0 ��[�i�e� O2ODOVO hOzO�O�O�O�O�O�O �O
__._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o[/& 8J\n���� !?����"�4�F��X�j��?[��1������������ q𩱬���Џ��� �%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A�S�e�w�L���Pӂ� ��ѿ�����+�=� O�a�sυϗϩϻ��τ��������#�-����j����	�12345678�f�h!B!+̺W���p�� �߷����������#� )᫿L�^�p���� �������� ��$�6� H�Z�l�}�;������ ������0BT�fx�����BH��/A Sew��������//��;�j%/O/a/s/�/�/�/ �/�/�/�/??'?9?0K?]?o?��D�y?�? �?�?�?�?�?OO1O COUOgOyO�O�O�O�O ���O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo�O;oMo_oqo �o�o�o�o�o�o�o %7I[m,o� �������!� 3�E�W�i�{�������Ïa������ׅ���0�B���"C� A}���   ���u2����} N��
���  	�a�2ޏşן���
�K7v��������1��3 4 5 6
�g�y��������� ӯ���	��-�?�Q�@c�u�������:�Pβ(Բڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�}���$SCR_GR�P 1C�|���~��t �±� {�	 ���� �Ҝҕ����}���G���������Q�������D�` D��@)���@���7��R-2000iB�/100P-IF/ 890��q媐�RB1P 67�8³
V10.'03 ����"�����������¶z���z�7�����������	��1�C�U�g�y�´?��H��������²E��BrLwDrR���3���g�c｡���ѺT�����FB���T�;[,��18����  �@��AE#+�B~;�Dq|��е�±��>��b�W�S���B����B�ff��  �����Au�� � ���@� � ?��c�#���F@ F�`N VMze���� ���/��G/02/D/V/h$B�v// �/�/�/�/?�/?:? %?^?I?�?m?�?(��: $����7�?{����?h+O²@DA�g1O���@1�kO� ȁG�12345��9A0�GHݏ�O´A ��6�E��r��@7���± _._@_NZQcXo_�_P_Ϳ�_�_��\Z�EL_DEFAULT  ��?��V��P?HOTSTR�]Q��QMIPOWE?RFL  z�j�1`WFDO�V �e�RRVENT �1D����"e� L!DUM_�EIP�_�h�j!AF_INE�P<�o´!FT�o�n��o!z�'6{���o[!RPC�_MAIN\>x�8J�nsVISw=yy���!TP�p�PU��id�?�!�
PMON_PR'OXY@��fe.�����Y��mfz�׏!RDM_SRV؏r�igƏ#�!R�Dd?��hh�o�!
pp�M���li^���!?RLSYNC����8���!RO�S�o.��4��S�!�
CE�MTCO�MT��fkB���!	�h�CONS���gl쎯�!h�WAS�RC�fmگ7�!�h�US��U��fn &���"���t���п ������=��a��W�RVICE_KL� ?%yk (%�SVCPRG1�hϰʚ�2�ϵϟ�3����ϟ�4 �ߟ�5�(�-ߟ�6P�Uߟ�7@x�}ߟ����߻�9������:��ߟ���� ����E����m��� ���B߽��j���� �������5�����]� ������3����[� ������������%�� ��M����u��#�� ��K����s������ m���Ϙ�8}�� �������/ �5/G/2/k/V/�/z/ �/�/�/�/�/?�/1? ?U?@?y?d?�?�?�? �?�?�?�?OO?O*O QOuO`O�O�O�O�O�O �O___;_&___J_ �_n_�_�_�_�_�_o�C_DEV ~yi�MC:	h�N�dGRP� 2Hye`��b�x 	� 
 U,k`�p�_`�`��`q�	o`pb �``�o�n
��d�a�o�j �d�e�k�gq-�a �a�o@�J}Ru� �g�a���i��{nd�   �Xp��`e`�d�  �`9a�Q�hJ� � ```(�xXs	`o�* �cB�j����g�a��ʅ ���g����B���� �aʏ ����i��LwhB�͟$���pXp�J`>`G?��� + `R`(���B�k�d&�Y��g�d@.��kB������o ��ޯ���(��L�^���fr���&��_`�`c+����jV`�����`@��"�� C�@ϛdj�2�D��yz� tϖ�����z}�τ�*����"C�"�	UXp�*`���`L���b"`�^�$�v�� �ߺ������u�� �v� O�6�s�Z���{��0�����"�v_`�с?`�ֱ�a���c|�d���$����h�Ρ ���d�����eƟ�� ��n�����c��n T�$���y� 6H/lS�w� ����� //D/ +/h/z/��/U/�/�/ �/�/�/?.??R?9? v?�?o?�?�?�?�?�? O�?*O�/O`OO�O kO}O�O�O�O�O�O_ �O8__\_n_U_�_y_�_�_�_�_CFd ��Ta�e6 2���>��>����R�����%'>В1>�����Z`������B.�S��nec�.<�����/m�	^�%fAZo�,��U���f߰C;F/mB��Z8B7!r�����Aҵ+B���BA�Y%�S103_PK�_TCOMUM3�5_R01�_s�#�Te:h`;a��~_�W�r��O���k�����O=�?�����u;a?!����Z�JAr!��@�����ߥ��,^}B��dC�?A����B�ES�k���A�	[~,��A�ä����V�Ü:A��e��S/�y%�
PRT46PI?CK1 N1�o�w�/Te<��e;����;t
�;��P�:��;.�.*;A�;}���zE��:A�j8�@x��W��X�+~����@�ݐA���B���V'=AӔh}��҃�AO#����]��E��A�r���	F�{�tS�ot�LTe�R6�;a<��䑿V��4`�<�0�uo���+{�~��\	���QA��0?�`��p�>R�Z}�������B�O�CKB�Bz�BMQ'�}�:MAG���A%��c�2@�@4H�O�JOGGI?NG K  �oI��TeUO�e>@�y�+߿}F����K^��g��;b:���K�j���A���@VrS���ߒ�>��ӎ��l��B����CC��Bf��;BBp}@E�[YA������\��I�A�?:??��#�5���Y�x`sr��?o�?����?��ſ��F��d
��T��W���wA����@X4PA߄A@�~����T�cH�B���~B(��<��C��`~���jA������t}���T����tO�6�PROC1��V�/�3�;�s�;���g;gӓ;����xG��V1�������:�A�@����A��@�Pv�����c�U�B�߆B(�n��;��C��wu>R9������?[�-���V��&��˯ݯ¿�3�:���H<�{B������z5_�>�Ѻ����~���Z��,pA����AX�A��#@_<BO�����cT�B����k��o��C� ��~Cz,A�`�j��]�I�����K���������p`r�[��V����n���E���������L����#A�<�A?�������?�T#�ٲ.��w� B8�?�B�|���uc�C]`J�CAA���p�F<��g��{AuI�?����sυ� ��l�HT�e��e?0��?�Rj@W1�>�В�q��5ʧ�������*BA�i�>K�A`���8�#���Î���yB�i,C��B?���B�r�;a���p�A��d���ޗ�9�����@]}+���	�P1 CON�VEYORl�V�l�:T���r��i��Q��?5+���7ڐ�g���?}.~����Ђ���A�~}���h�?*�+~��W�°�UB��nkB��r��:��k=��~����A��*�ߜB���=�"��i�yѤG�S�18�r_REAR�_UPPE;�CB,�Tl�83����@���@�B<�� <���F�@A7���������A���@�M�eA#�����R�#��1Y����LB�HC�����6X�A��o��~;�y@��U�������2�)�`|A���~�%�p50���_V2 f�CF6�'�A�|��<����Q���J1�r�<~����`�����A$p@�t�A"_{��"�s�*���B��1mC����5�A���~�T�����������js�Л�������H۶n�`;��m�<[{���ZlCA��~���$~�A�@ss?AJ����W �q˴B�2��s�U�5�cA����Ϟ���A��Fg��������]����>�pͤc���I�eCA;��2�YVZ��;��}Zl:����3���@tTAgW����*p/U�3�7\?�}�=p�^A���������\���X@Ygy������3�>�ɪ?��M�@�^���ɛ��?�Q�n�$Y����A��*�v�����]�RB����C��k�6��A�Ҵ~4�����I����Pp��(�&�K/]/CD;�w �{&�d�?��M�?�,������O�?G�����2�����A��W���	��/���YB���� ���6�&A�Ʉ�~J��A%����f~�i��\���#���?�7�A9�Ƌ����t���^��� ��A�Z�¿?�O��W~�@������QBt>��>�!�?�x�#��p���Jv�B��e��62��J�A����#��Aq����|��?���Mٺ�?�u�?1?�T!�Tl�B�e@dj��@
e��x����e�@�	���֖�~۸�I�t�A�4�P@����Q��?�:�#β��7��B����CAmB��a@N//�~� ����$�30O��G�y�V�?��V�G�50DR�O1��ϴYCTn���W�>^�T>�g�>���=���T=��;=��"��q�UmA�vNS@y���}ɿ�7+~���D@ǖ�A��SB����V�?A���~����AB����4��a&B�'b�H���	q1�q�P5�hRT�s~��F���,��? �>�:�X�:F�����h���N�An��?�Z}����ٿ6Β���C�<+^B��L8�b����>�0���~��z,@�ᒿ����(�?
��?r�G��FANUC_L�UB_J1_J2�_J3 �_��T�s*�.���	$�B�ӷ�����;��];���;�o�����{�A�?����}�(����n[���B΄�8���Fp:��mf^��jA�L g��R��q��0q`mDV��Ty��/�F�b�?����@qGC@���V?�z#?��B�oA��j����5A�V@��zE��ɂ��B���@��4A�1�B���f��A���Ξ�'��@���������'�qB+�����@oj�_�STz�A��E������}w�.Ƃ���[=�<��r�.��v�����A�Ʋ���p������7��������]�B����̐N¥�B�=��ϞVE�A��!X�HZM@��33�z�?�|d�O�O՟��zVߓ6 *�b��޿�n���U����Ꞿ���7>���w��m�L%A�z@����@^[C���J�g����¡� B��A$��Z­�Y�r��)^��mAr�J��$_��3��>�����C�G��3OUN�CE`߬�Tzz�+�V��`>� ��?��>���>��=����^�`����A�4+��3J���ȼ?����n���Ahx�A�mrC4���$�©�c�.�tX�A������6�D�OA��Q��yߎ$� waO����1��F��ť>��6?�y�>Գ�>�3v=���.�����z!A�8�οHbo��9<?������	Ag�)Al�,�CX?H�©�I��(!�c9�������5+SA��T���E[�m�����~���Vi�m=
�]=��>{���=��A<�P�Y^�$l�jp��@���������6Z?��?�B�H*A3-$�AջC���©
I­ȍ�^��jA���tz����A��f��=L�/�m�&� OT?�JW徭t�>3��A@I5��5�Zg�@ ��fo���p�A����Ay)�?���?����n���_�~\1B��:OB�����n��r�o���gaA�N<���7���� �@2�X��������� )TP��W�"ia�J�y�@������ɿV��@���oT@�����A��AA�����f�_A�n�����z4�B��B�1_���{vo���;A����{���'bvA�C���x������ *T�tݧ��qh,�G>�_Ѿ@���6�o=ք����HA�ja@>�P?K�h@�p?^��7�A�B����A@J����B�����0���P����V���%���2�t��JO?GGING �_���T�J��E>�n�<@	x]@8l��=ϱN�x�|��̆C9����1nA`@���B�?��>|,�r���w�^ �����6��&BAn�.���yA1�g����_@�xȿ��Y?,������3�T�~�å��`��¾�%��������F�ϳA��BN3�����A�a@��H�����>��־>B����!��0B�;B��"�d�eB
�'d^�p�@ �������"��-A\&����$�job38voK(�S^�bå�n�`�e��g������Žc��=�$�V�������lk@�i��@1����A�Z}?^���As���@H��º����	�C2���;�>R�����B@d�I>����A�@��m���@	�h]��#F���B���Bl�}���$��B9��~�?���4�A����A*��@V�rS������!�B����B�1��f^��³\Z�����A|����"����>�&F���^t`g���	�St|����	��=X? � ���'���?�@���^d@���k'A�ز�A5D���a��?x �n�v���Bc�B��-��)Bi�9�;n< @�u���%Q�r�.A,�� �Z��3�/�9%Swp������?��t���Nc@8�i�>�0�@ ��;n��JA⇿�@���X�������n�`������B�`~B�B����B�U*�;n,�������O���E@T@�Ͻ��&�����/�w�p
7W1H>mP�:�}�i?��=zb]>��~��bw���q��A��@�N?/��'<���'O�<�³��B��i�BB��G@4�BU���� �ۿ�	{�<���@��ҿ��!{wO��_STA�35 �O�I��\��>y�ؽp���?�s=v�l��O�`d�7���	�A��,@��6����;1��n���³�q�B�z�BB7����BT�@�W�J����$��\�>��@�?��V��K_�OBo�B��X���>y3������?��=���E>ғF�O�@����A�AQ@��]��P�԰W�_���³��B���eBAل�߬BTQ�W��)����`&}���4�M@��"��Ho��K _�/�M��YZ>�noU�x s?��=qz/>���"���P����?A��.@���(�������<B�ox�³���B���BA�{���BS�����ʟ�#�3��M��<{c�a�����o>��T20N1=b?o��F��ZE�>y��l��Q?����R������o���sA���@�Q�m1���4Pw6�³���B���BA�E��BS��g��T���ߞ�7k��b��7�Xou��Mq� å�l��Ǽ�?9jx�vL���(�8>��<��L�inA���_AP�?����K�B�;@,B����BA����+TBRn�W��%ga@a����r�G�{g�@�%*���ڛ��s7o�,��v����;|��;���;�[�:����:ݯ:A��;������As��@�>L���_��߾����@�IA�?#�B����T���A�T]�����APe<_�2�)S�Y��� �?h��QS�N�7%�D�/6�z��z��S���r�Ϳn�@���߽���g�:J��n-$�5�AϢ���h /������1?!��B�n¢[B����Cvc�W��3� @��@�� @������#9��<�.38DR�O��<�T&�����?b���%�)=a|��O�վz�
��T�aW��Qh0A�W�A"_{?԰�@~�߾_@c�¹!@B����B	n¡���@W�6s��!�����(��1��@aZ$������S198�0���'��k�@���@���@�i;�K^�.�_Y��ʧW�(���� �AW��3J�=`�>@�w�/�!����5�BYl�=��#²|��)��s��u��S���?�>��
�@��K��N	zj{���'���?�>��T?���>�9�:��a\������tW������~}AN��v�?*�@�h�/� �a�����BY��=��W?²z��)���s���*�>4���&?�l@�zP�!��ґ�2�������m?{8`>���h:����U�!����s�`������ANQ�#��?R�Z@�Q�� �N����BY�Q=��l�²q(�)�}Ʈ���&��>����(���G��9���1d����������?���S>�������$��y�>�����vA�Oja�Y�L?�8�#��MS����BZ%S=�{�G²e��)C�����!Q�s?K,�?����@hI9����8C�S105_GDR_�0�`�/#���c�!��8��R`/�!9}Zl���FV.>����V:A�*ҵ�<о�?�ů�� W����B�Z.=� �¿�h��)gFξ�4pƾA3��?��>��p��}+g��rC������w��,Cꏿ��8���݋!��h�����A�D���"���K��h��W���O��BZ�=�E=����)jf�{��Af]g���!?�����Y\/ �����w�:X @�0���5_�%�  ��Z.�A0o_���L�,����W�� SBW�1�=Ѥ�����)�nj����H?��a�?I�?�?�ʿg�n�1o�����w�!�(��B�9z5_9������ܑ7wQA��Ӑ����:R�>0 gW�����BX)��=������)�q�#^҃�=����+m�?7�}�?�[�>�`L��r41T����׉�@��_@Z��'>�9/==�Y��h�A� [AZ}>�0;/�W���CBX�|=�:�����)t��M�4P��?r�W�?WMuA?�/��/���ׅ�9�� ":J@ ��Q���/ <��} �jOAK=�����Z����>�Ơ?W�����QBX&C=��|���l�)v�"���^�-���s"�������_?�VO����S�p!69e�⻵K94�c}���}����rA�N���{h���>}Ǯ�ɰ��?=BX"�=��^��P�)y�?�����MA���0O>ǌy?�&Fc�詏SO���S�qY��{B�au-Ys���t��
VA�������˾���>X��OUg���=�BX �=�+��3;�{�.@����m�u���>���?4H�w>S_!�_����ׅ�}�9���gӓ� � �?1�`��E�wA�0R���>�oN~�"�����<''0�=�S}���)����]�@۱�Aww�z�z��_��_�_��,u�'�h�@��4H�?"��L�2G���?�޿��?�`q�l�gA�:�A�$!x?�L%@�fD3�. �����[B�cqB�9��mA���y?���Ay��2��¯���JO�{+T�,x嫐2C2#��½��̽�*����L�=]��<�_��A��rA��)jB �4�?�P@���@����4t�����B#���C�Ů�pM���6`�Ǯ>��A�(y�O�r�����^Q���F
z�o��gx��u����D���|m��wj<��=d��A�Y����f�A��?p@��Q�@��:��g�����B#��
C����ps�Y�6e�Ǯ5C�JA���G��ڿ\�����k��W�i�N�.��1I����2� ���, ����p�3o� ��v���o�@�?�����X�>��������(��@�钹qf�??�������A4��A5�o��k�p����o�o?Q���3M g���nub?]����1@)`Y>hT@��O���?�0��ɔB �{/AH���/�Ơ?"�������§�B���BQu���YBD-��p��^@��<�7�k���Qe���i���6��z	�%�41�� ���g�T6HVg��[~�y>���=�W����w_�X߄>P�.[�Ơ�s����A�J?�������7���	���I�A`Y�����;����C
[�i��@2D��E��?��A����m�zI�3�_PK_A�̼dT�6X��������-@j$���=@1�r@�%֞����Q,�^A�LA���,�f?��ێ���\��pB��2B�)�¿�S�%��� TA������s�>A?����O���������E�(g�@���>�c7�>�����T�?�?_�? �?��5D�A���@X4P����￪��/��)]���?B�M���k�Ԓ_���v?m��i���m	{�����@�Y�����RET_�HOME���h��THd�CV�W*����L>������Ⱦ<Hs�:�?�VrS��lk'A��t}A$ @-#�@���ێ-�¶˕�B���B���	A�"��S�e������A���TYF��؋V��}7�s�Ϭ}H�x�i���am����2�\��?�۹���X>����[�����r�B�{���Ap���$p/�J����<�B�eZ�N�������c���zg�8�A�9���c�A%jW�c��@�ޅ#�oDROPD�5 A�h�&TK'f��L�?�V������@9u>��r@��>?���)��ymA����@�N����dy��ێt����41B�yVB�89�FB�I��.�`�1��@����O��@NH����{�EO��E LFE��6p���,k?��k��=� ��?��?�sc.L����|OA��C�AS^��Cz��rz���jL��GB\�B���i�Bq�+7n�5��A������8��~�A0В翍�^;0�1 C?ONVEYO�t�LG{�)�	��@���j.�0��1��An��?�"�࿬B�@a��</��3�
��;A�d���{����q�xY����Cz,�f�����T��l�@!6��_�U_���G}�*?�A?�u�5__����x�A�_D<`�>K=�_�22��A�b��z�C��ydg�>�Q��zm��k���!@B&F�$a�ڊ������He�:2�H�Y���3�I�20`��P~�1N��Aw/��O��!�2��	(߮A��� ����M ic^���@��@���⼨
�@GY���-_e/w(e��p�?�1?��=�+a:>џ/�����9<A21\�=��翟����1�/2�����A��s ����� o[���9���j����2&i���*?<?�z%�#�z�@%�9l1�:����� �����AL���p�ǳ!�?2��N_A��� ��0��?�P�p����t���� �(>0
��=�E/�?�O{$2��� �"����P�:�X����tӣ����t�AT�W=L���2i�@k�)�sO2q�L��A�����B�����a�0מ�]���C�m�)O��=�@�Y��b���O��_`N���I#a:�ޮ�U@���[�!���� �A$��6?�?�����/���&ARA�<����1��~6� @�/&�@E[�Y�H��@�0�>�@�j�?L��H�8��]��	�2��@,�{�����ք�م�@�'Ӵ>l�K���o��AwA��:~��2C�~�7�@�"�g�Z�EA0b��;ظ����C/9��o�V�W5P�<��.�p��p0���o>}9 /���A�HY>����?��,����o��A#A�~�z��3r�~:τ@���7��f�]g�4���"Pp=<�De�_�X�0+IP�J�!�9�5_�� ?��!�.8�A�S&�;Q?��fD�3�eA��A�.���4���~>�@������	5¿������a�;!�<����n��Q
��I�4{y�Q�T�!��<����Β��AK�h�1�?�2�@o� ���DA&A��,���5��~A�@�t@S����ADxA�"���|��"�i?p�F+�)��V�|3���A��?�`��v���-���U9���������s����rAU�U�@�1X�?%��B��$@�K�A���B�_w�[?şA��Uw�P�A��[�������.A�� ?C�ӯ嫮�P��4TZ9.W5�x����座���s���HĿ�e�?�*w�X��u5A��X�@�_��տ ֿͨe�ޤ�O��ԡ�A��@�B��w�r��SAꈍS�;�yA���؀����鉿|d���

��6��_��/�TZRD_��p���r�~=�����ؾ����n?�������A����"����?]zE�����²�YBP��@C9rB�LB?�����"T`}�0�{%y�0����@�Y�c�6� �\�<TZ�|_�"e��;�"ٹd�� �o���R�Z��~}A��D!Ach���@ �? ABR�³�bB��=�Bߧ��ȍ'���?�'�@@��YI�Q1?�72=��MMOV`ҵ |P�0�TZ~'_��Ƨ�>���>�e����?�S��3J���mA���S@Kj@��� ?l@��������k�B����C8��B��ߎ@�wS����������c����gq�)�?�g�7�I�� *TZ��_�����>�5�>��Rr�m�Ľ�6����S������]A����@=ք@�!��?���n���IB��l�C8�Bů��?�F�wЀ�}����tz������?�������,TZ���W5;�!�@���?�J�?f���>���������+����?�$A���A`����A�@AZ�}Of����A��dB�]���w<�B���Β_|A�D��&�����LAA�U�S/:��o�ԑ���bTaB��W5=�,0=����=�g=��;='@�=&}��>�Ơs�T��APK_?��L��!���B��,�@���AѪ��B�*p�Sei�A���~i��?�������yA��x����38��E�������-$=��F=�=?�0= S8��Ѡ��bo��`/A�T�?���ވ���L%7���Y@�^4A�6��B���S�߃A�sQ�~%g�a=����,"�P����A�?�=�h�o��ʠ �2U����:g�ӓ:;��!=�������A~�o�A#x���{�����"5L����	�����AN+��ۋ�����C����>҃�׺����B�H��{ɣB_�G仟��C���a�2�k�!�=S�e��6�o�ٹ�=�� ꮿ��A�ۂA�������A;�H�� վ�����AN����ml���yC�~d�>�����i�[f~B �*��B^�Z�!/3("�m���O�/�V?�VY=�I������~2�A���AW������A�(��_���$G��AJ���܋����} C���>�ga�Ɩ�r�VvKB*�����]xA�Z���/�Cs-.5?&��UT�6��V���? ��=�?����_a3?E0��ecA�:����K@�)��9[?�t���AJ�����r����C�[R�?�0�K9����!B*�����A�廫?R�4S�//,8k9�`�?*>ICn��&�v��Z��>�ph�~�x����JA"����)X@�����!~6�� ��6uAQ���_1�����ef��,������(�A�nG�˯B`��O}ov_�9"M�FX�>�t2�>4ol��8����>�&���Ψ�����V�@����zB��@�/.�ʐ�_��;�A�QB���e����%CY>�����<��U�DD�B&F@���S_�e[!�Io8#O9�(� ��S>�0�<�3v���Q2>�"A���A|O�����r��@�yfޗ �S��AL����I:���a�C���~`¹�a����B(I�?�?&FA���'oe_�9"Qk?���>L4޿~���]p>��^���������x�@�#��h>p�@�;|�!b]��o��o�A�R7��������bCF�?��������!A�x���|AB_���o�4|��.-Tk�0?�K�?$y{�a~�����?��,��NH� 0��@C��x�X�@��
��0������{ASL�@��U� 7!C������H����I�F<����\=��@��];�Ə�!��$SERV_M?AIL  ᓡ������߄OU�TPUT����@߄RV 2I|�����  (w���x   W J����S��y̉߄SAVE�zb�T��0 2J+�� d 6E ee����
� >G�W ����?��W �G�%���W �G�r����U��������G�U-�����7GН� &T��*J��$�'��G���Es��`G�1"����
G�.��;r $�i����c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�Iπ[�m�ϑϣ�1��Y�Pn�a�FLT_C_URGRP�?������IDX  3�� 5�$�2�N��NUM���
��_DISFU�����ERR���?������o�TIP���Ӽ���ON  ��������SCH� 2K3��
2�'� �`��ԃ 2�4R�d�/�}��2� N����������+� �O�a�L���p����� ����������#� 5�G�tk����� ���(L7 p[����� �/!/4/?Qc �/��/�/��/�/�/  ??D?/?h?S?�?w? �?�?�?�?�?
O�?.O ;/=OPO[/m//�O�/ �O�OO_�O_<_'_ `_K_�_o_�_�_�_�_ �_o�_&ooJoWOYo lowO�O�O�o�O�o�o 5o"2XC|g �������� 	�B�-�f�sou����o �o�o��o��Q�>� )�N�t�_��������� ��˟���:�%�^� I�������������ӏ  ���$�6�m�Z�E�j� ��{�����ؿÿ���  ���V�A�z�eϞ� ������˯ݯ��� @�R߉�v�a߆߬ߗ� �߻�������<�'� 9�r�]�������� �������8�/�\�n� ���}����������� ��4XCU� y�������� �'�TK�x��� ����/�,// P/;/t/_/q/�/�/�/�/�/�??�$S�FLT_WAIL�IM  ���  ��;7TF?75REC�_GRP 2Lw����1r x�/�?�/�?�?��?/=ZN_CFG M�7w2:(6�D�2N�9�q,B�   Aa@D;� Bb@�  �B4RB2�156GTDSCH� 3O�5S3 �  �5�1�O�O��O�O�O�3 �4_+_=_O_a_s_�_�_�_��;0H7ELLBP�K��? '?o%RSRoo1ojo Uo�oyo�o�o�o�o�o �o0T?x�a�X1o%��Qcia�L����r2�dsra?��VHKw 1Q�K <� e���b׏���ޏ ��,�>�g�b�t����������Ο47�SOM�M R�_���FTOV_ENBi6� t5_�OW_R�EG_UI?�92IMIOFWDL
�AS�dEt�c1<���\o�c1OUTi6Dܶ�f8��ӯVA�L��r�_UNIT�;�
�t9LC�PIOw 2T�K�!� l�~�����ݟƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�4K7�`�r߄ߖ� �ߺ���������&��8�38@�SU 2UJ�\<�Q�\x��y��)����7��  ���������+�� ��[�m��������N�LERR 2V�IH�� ��_�� !3EWi{�� �����/ ASew���� ���//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o?��?�?�?�?G�Y�TR�Y`�J�=�MImSA2WJ� ��?�����AO/H^Ѹ���
�t~��0C�O O��O�O�O�O��_IR�D_MAP  �n�YOkA�PMB_HDDN 2Xn� }���S]I_ [_�__�_�_�_�_�_��_m+QON_AL�IAS ?e��( he��[omoo�o �jIo�o�o�o�o�o .@Rd��� ��{���*�<� �`�r�����A���̏ ޏ�����&�8�J�\� n��������ȟڟ�� ���"�4�F��j�|� ����K�į֯���� ��0�B�T�f�x�#��� ����ҿ俏���,� >��O�tφϘϪ�U� ����������:�L� ^�p߂�-ߦ߸����� �ߙ��$�6�H���l� ~����_������� � ���D�V�h�z��� 7������������� .@R��v��� �i��*� N`r��A�� ���/&/8/J/\/ /�/�/�/�/�/s/�/ �/?"?4?�/X?j?|? �?9?�?�?�?�?�?�? O0OBOTOfOO�O�O �O�O�O}O�O__,_ >_�Ob_t_�_�_C_�_ �_�_�_o�_(o:oLo�^opoc�$SMO�N_DEFPRO ����a� *SYSTEM*`�49�dRECA�LL ?}�i ( �}"o�o�o1C �ohz� ���U��
�� .�@��d�v������� ��Q�����*�<� Ϗ`�r���������M� ޟ���&�8�˟\� n���������I�گ� ���"�4�ǯE�j�|� ������ĿW����� �0�B�տf�xϊϜ� ����S�������,� >���b�t߆ߘߪ߼� O�������(�:��� ^�p�����K��� �� ��$�6���Z�l� ~�������G�������  2D��hz� ���U��
 .@�dv��� �Q��//*/</ �`/r/�/�/�/�/M/ �/�/??&?8?�/\? n?�?�?�?�?I?�?�? �?O"O4O�?EOjO|O �O�O�O�OWO�O�O_ _0_B_�Of_x_�_�_ �_�_S_�_�_oo,o >o�_boto�o�o�o�o Oo�o�o(:�o ^p����K� � ��$�6��Z�l� ~�������G�ŏ��� � �2�D�׏h�z��� ����U����
�� .�@�ӟd�v����������K��$SNPX�_ASG 2Y�����_�  0R�%X���R�?�զPAR�AM Z�^� �	��PK�eR�K�`��נ�OFT_KB_CFG  K��ԣ�OPIN_SIMW  �[����ǿٿ�נPOTT�SKINFO 1][� ��� &�8�J�\�nπϒϤ� �����������"�4��F�X�j�נRVQS�TP_DSB���[���̫SR \�� � & �STYLE103�_TC 4_J5w_J6�� Ѧ�TOP_ON_ERR  �֎��PTN ��>�A�RI�NG_PRM� �נVCNT_G�P 2]�]��x 	[���K���౼d��� +��,���+ˬVDm�RP' 1^4�^���� ���0�B�T�f����� ������������ ,SPbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?k?h?z? �?�?�?�?�?�?�?
O 1O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \o�o�o�o�o�o�o�o �o�o"IFXj |������� ��0�B�T�f�x��� ����Տҏ����� ,�>�P�b�t�������༟Ο�����PRG�_COUNT��q�>ᑵ�ENBS���MC���P�_UP�D 1_��T  
�O�������� ����/�*�<�N�w� r���������̿޿� ��&�O�J�\�nϗ� �Ϥ϶���������'� "�4�F�o�j�|ߎ߷� ������������G� B�T�f������� ��������,�>�g� b�t������������� ��?:L^� ������� $6_Zl~� ������/7/�2/D/�_INFO� 1`��n� ��g/�/�/��/�-<3��V%����'�%�T����FB��T��;[,�18�k���YSDE�BUG(����] d�q�90SP_PAS�S(�B?K;LO�G a�&s�z] �1�^��] �d/  �m�]!
MC:\w4x3-;z0o_MPC}? �4x�2O�<UD1�5�2k.�3SAV ab�=�!�1 J'H�SV-;TEM_T�IME 1c�7�t� 0 �C�]"��V&�v�V',��C`Rv�T1SVGUNS���)�'q���@AS�K_OPTION�(���m�u��A_D�IZ0D�UBCCF�G e��R
J�" O]Z`{_�/�_ �_�_�_�_o�_1oo Uo@oyodovo�o�o�o �o�o�o+Q< u`������V$�|��@�R�� /���s�����Џފ�� �Pŀ����B�0� f�T���x�������� ҟ���,��P�>�`� ��t�����ί���� ���L�2��`�r� ������2�ؿƿ�� ��2�D�V�$�z�hϞ� ���ϰ��������
� @�.�d�R߈�vߘ߾� ���������*��:� <�N��r��^����� ������8�&�H�n� \��������������� ��"24F|j ������� B0fT�x� ����/�� /2/ P/b/t/��/�/�/�/ �/�/??�/:?(?^? L?�?p?�?�?�?�?�?  O�?$OOHO6OXO~O lO�O�O�O�O�O�O�O �O_D_2_h_/�_�_ �_�_�_R_�_�_o.o oRodovoDo�o�o�o �o�o�o�o�o<* `N�r���� ���&��J�8�Z� \�n�����ȏ~_��� �"�4���X�F�h��� |���ğ֟������ �B�0�R�T�f����� �����ү����>� ,�b�P���t������� ��ο��(�ޏ@�R� pςϔ�ϸϦ����� ���$�6��Z�H�~� lߢߐ߲ߴ�������  ��D�2�h�V�x�� ���������
���� �.�d�R���>Ϡ��� ������r�(N�<r\� �$TB�CSG_GRP �2f\��  �� 
 ?�  ��� ���K5o���h�d׼^�?�	 �HD)��a��� �A��8���333"���B ��
/.H�>/�-Csx^ �%�CA�t/D�/�*Y��%�' �/?�*L��46�/R?^8@�_��5�?b? t?�?�?�?�?
O'O6K��%� �  	�V3.00�	�rb1p6C	�*r@jD�6CA-/ O?fff�A� x� ��I �@�M�O { i���CM?��OT�JCFG j\�T@[+�,R�B_WX�W_}_�Ze �_ �_�_�_�_�_�_oo Ao,o>owobo�o�o�o �o�o�o�o=( aL�p���� ���'�9����D� V�h��������я�� ������=�O�a�s� .���������˟� |�X&�(�:�p�^� ��������ܯʯ��  �6�$�Z�H�~�l��� ����ؿƿ��� �� D�2�T�z�hϞό��� �������Ϩ��@�.� d�R߈�v߬ߚ߼��� �������*�`�N� �����t������ ����&�\�J���n� ��������������" F4jXz|� �����0 @f�~��L� ����,//P/>/ t/�/�/�/h/�/�/�/ �/?(?:?L??\?�? p?�?�?�?�?�?�?�?  OOHO6OlOZO�O~O �O�O�O�O�O_�O2_  _V_D_f_h_z_�_�_ �_�_�_
o�"o4o�_ �_vodo�o�o�o�o�o �o�o*<�oLr `������� ��8�&�H�n�\��� ������ڏȏ���� 4�"�X�F�|�j����� ��֟ğ�����B� 0�R�T�f���o��Ư د������>�,�b� P���t�����ο࿞� ��(��8�^�pς� <�NϸϦ����� ��� $��4�Z�H�~�lߢ� ���ߴ������� �� D�2�h�V��z���� ������
���.�@�� X�j��&��������� ����*N`r 0B����� &�J8Z\n ������/�  /F/4/j/X/�/|/�/ �/�/�/�/?�/0?? T?B?x?f?�?�?�?�? L�~��?O�?�?,O>O tObO�O�O�O�O�O�O __�O:_(_J_L_^_ �_�_�_�_�_�_�_o  o6o$oFoHoZo�o~o �o�o�o�o�o�o2  VDzh��� �����
�@�.� d�v� O������\�� Џ����*�`�N� ��������x�ޟ̟�8�&��  L�P�� P�d�P��$�TBJOP_GR�P 2k���  ?��P�	|���m���� �� X��X��� ���, ��,XP� �@L���	 �D�)� �C2
�C랔P����Ù�$��%�7�;w{ �?L���A�b�p�s�~� ���4���ȵ<I��T��ư�BHb���j�ώ�����333�D�űA�S�;�]���i�B ����  �C�ƒ��/C�p���sV��������<+CA৬�}�d��-߰φ��?Yưe�a�s�;'����Y��V��� ����2�Dߦ�Y������<oܜޥ�F� ��a�X�ǀ�j�x�� ���l�������6� g�B������������d���ԇP�e���	V3.00���rb1i�	*�B ��K�P�A��[
� F�` p��0 F�  G �� G� G�� G$ G7�� GR� Gv� G�� G��� �� G�� �G�$ H
� H@ H.�k�� F;� FZ� Fz  F�� ?�� F����Gb� G�����P Gq H�� H(� HK � Ht� �| =u=\)��)xL����Z�@
RP�V���o��CPPACTSW�  ���IR �n��� C����SPEED �o� �/L������_CFG #p�O��P���P��_CUR_�ID頵�\`#E�XT_ENB  �L%x%`#HIST_BU 2q���dt��1'�7��(=�(C�(I�(O��(U�([�(a�(g��(m�(s�(y�(��(��(��(��(���(��(��(��(���(��(��(��(Ǫ�(��(��(��(ߪ�(��(��(��(���(�%(	(�(((!('*(-(3(9(̱*%E(K(Q(��&](c(i(o*(u({(�(W���(�(�(U�(�(�(�(U�(�(�(�(U�(�(�(�(U�(�(�(�(�M��chch�chchch#ch)�ch/ch5ch;chA�chGchMchSchY�ch_�(�(�(��(�(%�(+�_MAX_ANTm/� �`#SPD,#rtp-L���B:�BVaM���wNU�`�P�t)
�wOUT7 2s��
 YS) H�S%B�T���x����� ����ҏ���'��,�x>�P��ZERO�p��,w�ESTPAR`
p��^B|�HR��ABLE 1t���J/�U(Jh�ng  h�O�W�h�vG� h�zgI'�rh�h��G����RDI���q�֟�����0���O ������ί������S���s@��G ���$���0G!���O�k���PjA��3��W���O�na����O������0C$��O�3�1�C�U�g�J� K� R���@.q���"Y$�`�Dư����������  �2�D�V�h�zߌߞ� ����������
��.�@�R�d�v���N%� -����МN�K� ]�o���-�?�Q�c�u���B����� �
jA�@����,"�u�Z���IMEBF_TT��S��)��VE���G!z��R 1v�{� 8�9�r� ������  �	PRT02_2�74��]Dl (� �hzI9� ������� 1CUgy�� ��
/��	//-/�?/��T/f/@.GIN�/�/@/R/�/�/ �/
??W�Z�8?J?�?�n?�?�<nd�?�?�:��nb�?�?�:�� O&O�?�?\Oqr0��@�uspMI_�CHA� �� �u ~�CDBGLVL����v�CETHER_AD ?��Pm��0&P:e)P�4:3b:48:34 &_5oO3�:_e7TR$� !�z�!|T�_�y�@SN�MASKX�s#P_255.�U0kC��_�_�_nuOOLOFS_DI
p�����ORQCTRL w�y���so9�Tgo�o�o�o�o�o�o ,>Pbt� ����|fo������PDRAM��x6Tjd9����`� r���������̏ޏ��@��#���5��BD �5�K�)�E_DE�TAI�H=jPGL�_CONFIG �~����/�cell/$CID$/grp1#�@��ӟ���	�9�O_ 4�F�X�j�|������ į֯������0�B� T�f�x����+���ҿ ����ϩ�>�P�b� tφϘ�'ϼ������� �ߥϷ�L�^�p߂��ߦ���};����� ��$�6�p��^�=� :ߓ���������4� �#�5�G�Y�k���� �������������� 1CUgy�� �����-? Qcu���� ��/�)/;/M/_/ q/�//�/�/�/�/�/ ??�/7?I?[?m?? �? ?�?�?�?�?�?O �?3OEOWOiO{O�O�O����User� View ��}�}1234567890�O�O�O__�*_2T ��~�����NDeST?�]�B4  ^Q���I2�I/O�_�_�_��_�_�_eRo:��I3 w_<oNo`oro�o�o�_ �on_P-o�o( :L�oml5�o� �����]�n6�X�j�|��������ӏn7G���0�@B�T�f�ŏ��n8�� ��ҟ�����y�;��A� lCamera�J����@������ȯگ��Es� ��(��OB�T�f�x������y  Z�vYo� ����"�4�F��j� |ώ�ٿ�����������3��Z�*i��X�j� |ߎߠ߲�Y������� E��0�B�T�f�x�� 1��i���������� ���B�T�f������ ����������1׸�}� 2DVhz�3�� ���
.@ R��[�F����� ����/,/>/� b/t/�/�/�/�/c1� ��S/??,?>?P?b? 	/�?�?�?�/�?�?�? OO(O�/1׮��?tO �O�O�O�O�Ou?�O_ _aO:_L_^_p_�_�_;OMG9 _�_�_�_o o/o�O@oeowo_�o��o�o�o�o�o��	\�0�oBTfx� �Co����o�� ,�>�P�b�	a�c� ���͏ߏ���� 9�K�]����������� ɟ۟��\�ϻr�'�9� K�]�o���(�����ɯ �����#�5�G�� (u;�ޯ������ɿۿ ���#�5π�Y�k� }Ϗϡϳ�Z�l���J� ���#�5�G�Y� �}� �ߡ������������ ���l���k�}�� �����l������X� 1�C�U�g�y���2�l� "�������1 ��Ugy�����������   ��&8J\n�������   �D4�EJ!�d��?���B��D�P�?���E��@������7`ó=�����8�2���!Dol�@2��B��J!�@��kJ/\$
��A��3Aǒ`�R)Dz` R2Ae.�A�������~�Ğ�N�DeST@)<��A�h�B����Qév��̾��DM�@-��$A��B�!��Q��x����fD�]�@?�AW��%�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_�L_^_�  
��(�  �( 	 n_�_�_�_�_�_ �_o�_ o"o4ojoXoЎo|o�oxZ�
 �F�o	�?Q cu�����o�� �.��/�A�S�e� ��������я��� ��+�r�O�a�s��� ������͟ߟ�8�J� '�9�K���o������� ��ɯ�����X�5� G�Y�k�}���֯��ſ ׿�����1�C�U� �����ϝϯ������� ��	��-�t�Q�c�u� �ϙ߽߫�������:� �)�;��_�q��� ��� ������Z� 7�I�[�m������� ���� ���!3E W��{������ ��dvSe w������� </+/=/�a/s/�/ �/�/�//�/�/?J/ '?9?K?]?o?�?�/�`@ �2�?�?�?�3��7�P��+fr�h:\tpgl\�robots\r�2000ibE_�100pif.xml�?:OLO^OpO�O��O�O�O�O�O�&�� �O__/_A_S_e_w_ �_�_�_�_�_�O�_o o+o=oOoaoso�o�o �o�o�o�_�o' 9K]o���� ��o���#�5�G� Y�k�}�������ŏ� ֏����1�C�U�g� y���������؏ҟ�� 	��-�?�Q�c�u��� ������ԟί��� )�;�M�_�q�������蹿˾�8#1 ��?�088�?�˻
�˿�(�*�<� ^ψ�rϔϾϨ����� �� �*��6�`�J�l���ߴ��$TPGL�_OUTPUT ���!�!� �D PBC��+E(ZN?��+AR9D����!C����y?E	�&�@Qa´  ����%�1�C� U�g�y�������� ����	��-�?�Q�c��u�������23�45678901 �����������"���noselec�t*�!���A� )������d�Q����"|�vHB�!�P WD��EZ��Q�%���� hh0B���"�[� �.B�� ����� ��)BT fx�",}�� ���/��C/U/ g/y/�/�/5/�/�/�/ �/	??�/)?Q?c?u? �?�?1?C?�?�?�?O O)O�?7O_OqO�O�O �O?O�O�O�O__%_ �O�O[_m__�_�_�_ M_�_�_�_o!o3o�_ Aoio{o�o�o�oIo[o �o�o/A�oO@w����'}鱀���%�7�I�Z�@��~����� ( 	 ��ŏ���׏ ���1��A�C�U��� y�����ӟ������ -��Q�?�u�c������������������ ���M�_�;����� q���ɿ��8��Ϧ� (�:��^�p�ڿ|Ϧ� H϶��Ϻ����$ߎ� H�Z���~ߐ�nߴ��� 0����ߞ���2�D�"� h�z��ߞ��R����� ��
�����R�d�� ����x�����:��� ��*<Lr���� ��\���& �J\�l�p� �2D�/�4/F/ $/j/|/��/�/T/�/ �/�/�/?0?�/T?f? ?�?�?z?�?�?<?�? O�?�?>OPO.OtO�O �?�O�O^O�O�O�O_ (_�O_^_p__�_�_��_�_�_�R�$TP�OFF_LIM �3�h�/���h��RN_SV�P � a�jP_M�ON �+��dh�h�2a��QS�TRTCHK Ƀ+�f�bVT?COMPAT"h�a�fVWVAR �Bm�h&d R�o �oh�Ub�Q�_DEFPROG� %qj%ST�YLE103_T�C�o�j_DISP�LAY`qnrIN�ST_MSK  �i| SzINU�SER�oYtLCK��|r{QUICKM�EN�YtSCRE��p+��btpscYt�q	��b��_#�ST�jiR�ACE_CFG ��Bi�d�`	��d
?�j�HNL 2�qi����k �bԏ���
���.�@�R�l�ITEM� 2��� �%�$1234567�890����  =�<��şןߓ  !���`��2��c ��S���w���ퟟ�� #��G��k��=�ï ��ůׯ���u��˿ ��g�'ϋ�����)� ӿϥϷ����?�Q� c���5ߙ�Y�k���w� �����)���M��� ��5���߂��ߝ�� ������I���m��� ���a��������!� 3�E�����{�;M�� Y������/� e��d� ���;+=Oi s��C/i/{/��/ //'/�/K/�/?/? �/;?�/�/�/_?�?? �?�?G?�?k?}?FO�? aO�?�O�O�?�OOqO �OUO_yO%_K_]_�O i_�O�O	_�_-_�_�_ ou_5o�_�_�_AoYo �_�o�o)o�oMo_o( �oC�ogy�o�(�h�St��z��z��  ]��zq ��8�/y
 E��k�R����UD1�:\�����qR_�GRP 1���� 	 @�p ������=�+�a�O��q�����[�����x���ϕ?�  �� ���1��U�C�y�g� ������ӯ������`	�?�-�O�u�	�u������sSCB 2��{ ���� ��/�A�S�e�w��|�V_CONFIG� ��}�� ��s�֟�ϑ�OUT?PUT ��y������+�=�O� a�s߅ߗߩ߻����������q�Regu�lar Opti�on\R798 �: DRAM F�ile Storage�U�g�y�����������	�� �-�?�Q�c�u����� ������������ 0BTfx��� ����,> Pbt����� ��/(/:/L/^/ p/�/�/�/�/�/�/�/  ?/#/6?H?Z?l?~? �?�?�?�?�?�?�?O ?2ODOVOhOzO�O�O �O�O�O�O�O
_O._ @_R_d_v_�_�_�_�_ �_�_�_o_)_<oNo `oro�o�o�o�o�o�o �o��	����V hz������ �
��.�!oR�d�v� ��������Џ��� �*�;�N�`�r����� ����̟ޟ���&� 8�I�\�n��������� ȯگ����"�4�E� X�j�|�������Ŀֿ �����0�A�T�f� xϊϜϮ��������� ��,�>�O�b�t߆� �ߪ߼��������� (�:�K�^�p���� �������� ��$�6� G�Z�l�~��������� ������ 2DU� hz��������
.@#y���`r\K��@v  Regul�ar Optio�n\R798 :� DRAM Fi�le Storage��//)/;/ M/_/q/�/�/�/�� ��/??%?7?I?[? m??�?�?T�?�?�? �?O!O3OEOWOiO{O �O�O�?�O�O�O�O_ _/_A_S_e_w_�_�_ �_�O�_�_�_oo+o =oOoaoso�o�o�o�_ �o�o�o'9K ]o����o�� ���#�5�G�Y�k� }��������׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;��M�_�q�����������$TX_SCRE�EN 1�t�\�}P�rodHome.stm��
��.�@��Rϩ	PROD� HOMEY�}��YϚϬϾ������� ��~�+�=�O�a�s߅� �ϩ� ����������'�߰�http�://192.168.1.54I�������.�ATI TC����� *�<�N�`�;������ ��������g���8 J\n��	�- ���"4���/wizinst�������a��Wizard �Top Menu���UALRM_M�SG ?ڹ� ��  INV�ALID ARG�UMENT RE�CEIVEDŢ�$%DECISI�ON CODu��WAITING� FOR MAINTENANCu��Tip Dr�esser 1 �Disconne�ct Off@ ~�+Jammed����( G1 Cur�rent�o L�ow� � d�#(�s) Not i?n Auto}'�#1 Motor�"Start�!?4�opp2STEPPER NO3!�SET��Wa�tersav�"U�nable� R�eset`<2p>��+Phasev� ssǠ� "8��!Acnowle�dged WC1��?�:2�4�&2�-	�+2�+� J G2
�.	"82?�:mK;3P�;2�;' @L����AWTR 1:� WATI4OFF��M2�O�BEF�$4� Dump�3d/vanc�!"6+Y�Retrac1Y�"7N@._AXmXWW!8G�3n_@Y�XWWDbX4�_ 
BW�XWW�O��Q��-�P�+N�+3�+�m@L3PO"83nO �F�o4:�;3�;�P`D�&�P�+�+4�+��RG�*4�.�94F�o �b4:�<4�;� @Check� �%�SPin�  �K�d�sEqual{iz� Faul0� ��0$5� �%H�ighš� o�Cap Cha�nge ERROUR����0� l'���wyeP0 �Cou� Q�  �� Find�h�ŢP�2�Dn����55�3�����c �d�P� �!Q�e\�Search� Sens0Q�u6 @E��of
��~Q��ctOk1�Trj0ln���0�Anti Cra�s0�Ǡ� iR7Visz2rv�)Ǡ��0�����������0ß��� `㟽�/ @�¸��"�`������h ���`�2����0Key Sw�it�L1�!UTO�:���0Gun/�Backu1P�AP�հ2�� o2�xR �"�off det|� ���54$��s n�#the �c0ri�0  
�VAB�H�remoڏ�/mal�0  ��.fAdapt.z1iv�;P'��k�piz�OT�D Verifi�cation����0C�same a�s+�ach�"�$��2��2P�og�ram 0DIS�P_SEQ ErGror�0�2�� �r2�!@�2�� b��2�\�0��2�KDE �ϴ� `��2�̀ �ϒ2�G��2��`�2��$ �2��`�2�� �2��~ ߒ�pd��2�?��2�0��s�A�2�9� �2�#CSb�2�9�`�2�� ���2���@�2����2�tj99�2��""�2�9H �2��iob�2�9�`�2�os��t�Ia��2����2�F���2�r%1"2�LCIMB2�� 2� �2���2����2��0���2����2���2��PA2�!8A��2����\c�2��`2�A� 2 /2�f�2��`/���2�*@��/2�	u�/2�9 �?�	�/�2�q����2��\j�?2�5@?2��C ��?� ?2�� O�2�� ?�o��2�;�@/2� �O2��$�/�O2���?2�ɩ�/2�E _2��9�B_2�1Db_4�� O2�2  �_2���EF�_�Y9�_���RoT�R6"o2��$�_2�]@_2�I�O2�I6�o2���2���o�2�� _R�ao2�jL!VB��o2��@2�!`�or��2����@�s ���A�2��@���intShopN��@IF��2��䣏3�P�����d ��2�
du�2�\sfd"�2����B�r2�#�����_C���2�٠��2�?!ß3��Is�������w ����v@����`����s~܂�2�$"��"2�� �ï3�.����� Q@�$UAL�RM�V  ����0��� �  &D�C�G�L�O�t�z�&&z������Ŀֿ���"�ECF�G �0�.@�  ���= -��   BȚQ�� 
 !�� �� �A �SmZ��D�)Tj;�!�� ��A���T�P�tΔ��T�E�\��S�m���Sm����&Sm)����	 Sm*�~���Sm/=߿�SmA�	�G_RP 2���0�=�!�	 ��X�"���?�����`������6+�Z$U�I_BBL_NO�TE ��T?��l�R1��Q��DEFP�ROG ?%0�� (%	PRT11PICKm��X��7_R01����c� 6�!�Z�E�~�i������������z�INU�SER  �����_MENHI�ST 1��]�(~� ��'/�SOFTPART�/GENLINK�?current�=menupag�e,37,�01�_TC��35�,17A�������y����,74���Ѡ��EYOR��8J\n���,7�� ��2�N�V1���y/<���edit����50�3�4AS`e���46��� TE��,44pw��� �(�&��93#(3�P/b/t/w0/�+��	C��� E/�/�/�/�~2�/�/�&_V2��B!49?a?s?�? ��|Qw���?�?�?�? �?O|�?7OIO[OmO O�O O�O�O�O�O�O _�O3_E_W_i_{_�_ _._�_�_�_�_oo �_AoSoeowo�o�o*o �o�o�o�o�o�o Oas����?� ����'�9�<]� o���������F�ۏ� ���#�5�ďY�k�}� ������şT����� �1�C�ҟg�y����� ����P����	��-� ?�Q��u��������� Ͽ����)�;�M� _�b��ϕϧϹ����� l���%�7�I�[��� ߑߣߵ�������z� �!�3�E�W�i��ߍ� ���������v��� /�A�S�e�w������ ��������࿎�+= Oas������ ���'9K] o�"���� �/�5/G/Y/k/}/ �//�/�/�/�/�/? �/�/C?U?g?y?�?�? ,?�?�?�?�?	OO
��$UI_PAN�EDATA 1�����KA�  	�}�/frh/cgt�p/doubde�v1.stm x�.hr@FOC_prim'O�O�O�O�N#)O�O�3}�O_`,_>_P_b_t_ )v_ �_�_�_�_�_�_�_o �_<oNo5oroYo�o�o��o�o�6�� �   ! ���$R]O2pBg�.shtzBduaAl�o4FX�o��V_Fitree pB������o)� ;�"�_�F�����|��� ��ݏ�֏���7�I��0�m��n�`� KA_����џ���� Z�+��OO�a�s����� ���ͯ߯Ư��'� 9� �]�D���h�����@��ۿ¿����c N@ ,�MCH�M�_�qσϕ� ������>�����%� 7�I߰�m��fߣߊ� ����������!��E� W�>�{�b���$�6� ������/�A���e� �ω������������� \� =$asZ �~����� 'K������ ���.�/��5/ G/Y/k/}/�/��/�/ �/�/�/?�/1?C?*? g?N?�?�?�?�?�?�? Xj(/-O?OQOcOuO �O�?�O/�O�O�O_ _)_�OM___F_�_j_ �_�_�_�_�_o�_%o 7oo[oBoo�oOO �o�o�o�o!toE �Oi{����� <����A�S�:� w�^�������я���� ��+��o�j�6�o� ��������ɟ)]�� auݟ�,�>�P�b�t� ۟����������ٯ ���:�L�3�p�W��������ʿ[x�c�k�$�UI_POSTY�PE  �e� 	 ֿ�-���QUICKM_EN  ���0���RESTOR�E 1��e  ���Bcr�ϴâ�crm�� ����1�C���g�y� �ߝ߯�R�������	� ���(�:�L�߇�� �����r�����)� ;�M���q��������� d�������\�%7I [m����� |�!3E��� dv������ /�//A/S/e/w// �/�/�/�/�/��/? ?�/O?a?s?�?�?:? �?�?�?�?OO�?9O�KO]OoO�O;�SCR�EK�?P��u1sc��u2��D3�D4�D5�D6ʼD7�D8�A��UScER�@�O�Dks�C�T3T4T5T6�T7T8Q��ND�O_CFG ���F�E���PDAT�E Y�?None L���@�_INFO 1�2�e�P\�0%�O�_ [x�_�_�_o1ooUo goJo�ono�o�o�o�o��o�o4̞QOFF�SET �P� (C��*Ol~�� ������X� _�V�h�������ˏ ԏ�0�`�2�
!�V��4xUFRAME � DnV�QRTOL_ABRTz��8s��ENB����G�RP 1���\�?Cz  A��� sQ���%�7�I�[��m���J�U��sQ��MSK  ���RvQڎ�Nw�%�Z%	�PRT50_R0y1]�5�VCCM_R��f]�MRג2���ĐF�vR&@	�tPr~XC5G6 *q�{���sT֢��5&@sQA@�}�pq��� E�ǸѿH��1��^�,�Y�ʵk�A��$BEϖ�$B B��ͱ�$A��=� ��������	�B�-� f�Q�cߜ���}��߽������,�>��ISIONTMOU�����mU�U�����/��0��� FR:\�W�\PA\C� ��� MC��L�OG��   U�D1��EX��$A'� B@ ��
����(���,�P��C �  =�	 1- n?6  -��F��E,b�챝�=�S�ͦ�D����TRAIN��f��$A{�
&@dQ�9��@� (�Ѧ�"�� "0BTfx�� �����O�-_��RE��ޙd�^�LEXE��@��sQ1-eE�VMPHASE  �U�sS���RTD_�FILTER 2]�@� �2�Ⱦ� //1/C/U/g/y/�/ �/�/-���/�/??�(?:?L?^?p?�?�SoHIFT��1�@�/
 <�%��?h����?�?O�?O PO'O9O�O]OoO�O�O��O�O_�O�O:__�	LIVE/SN�APsvsflsiv�L_�W�� DpUiPoRmenu�_�_$_�_�_�R�5��ޚ	�X�_Loh㫲�� ~�@���A� B8��������ab��cV�:�@u�=��iP��(��1�MO����|���$WAITDINGENDb觨tO�����!w`�7SKyT�IM����v|G �}*�{J�zi�z<�xRELE���� t]�ȓ�s_AC�TbPJ��w_�� ���  NTR�IZONSo�o�R�DISiP���$X�S��ޛ��S����_$ZABCד�i' ,����2ӏ�WZIPc�i���ȟڟ|�MPCF�_G 1�� a0�[�"��MPB�1��ġ�$���z��8<o����j�ۯ��?�߫��߯ɯ :���a�#��������f�����ɿ߿�ˈ<����������Y�LIND���� l�� ,(  *xω��uϲϙ��Ͻ� ����0� r�S���w�^�p߭��� ������8��ߚ�O� 6�s�Z��ߩ��{�H�s2���� �� ��'���?�*�c�h�h���h����A�F��SPHERE 2�X�����]��� C���y�� N4��	�b? Q���������(//)/<�ZZi� �U�