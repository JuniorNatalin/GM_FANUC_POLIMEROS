��   u��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����UI_CONFI�G_T  �� A$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA}T��$TOP>�_IDXCMEM�_LIMIR$�DBGLVL�P�OPUP_MAS�K�zA  �$DUMMY62��ODE�
3CF�OCA �4CP�S)C��g H�AN� � TIM�EOU�PIPE�SIZE � M�WIN�PANEwMAP�  � � FAVB ?� �
$HL�_DI�Q?� qELEMZ�UR� l� �Ss�$HMI��RO+\W A_DONLY� ��TOUCH�PR�OOMMO#?=$�ALAR< �?FILVEW�	ENB=%%fC �1"USER:)F�CTN:)WI�:� I* _ED�l"�V!_TITL� �1"COORDF^<#LOCK6%�$�F%�!b"EBFOR �? �"e&
�"�%F�!BA�!j ?�"�BG�%�!jINS�R$IO}7P}M�X_PKT�"�IHELP� ME�R�BLNKC=E�NAB�!? SIPMANUA�L4"="�BEEY?$��=&q!EDy#M0I8P0q!�JWD�D7��DSB�� GT�B9I�:J�; k�&USTOM0� t $} RT�_SPID�,DC�4D*PAG� ?~^DEVICEPIoSCREuEF���IGN�@$FL;AG�@�&��1  h 	$P�WD_ACCES� E �8��C��!�%)$LABE�� $Tz jp�@�3�B�	�&�USRVI 1  < `�B*�B���APRI�mx� t1RPTRIP�"m�$$CLA�@? ���sQ��eR��RhP\ SI��qW  ϶:�$'2 �6|@��R	 �,��?�����Q�P�R�T�Qr�����P�@�?�^��
 ��)/SOFTP.@�/GEN�1?cu�rrent=me�nupage,381,10oko}ȍo���(1oCn952,1�o�o $��  �nCURRENT=>QA�ol@~��1CUu8_ ���)��a0o�oTb4-�{�����.���Տ �����/���S�e� w�������<�џ��� ��+���=�a�s��� ������J�߯����'�9��� /TPTX��zQ���g�y��P sO����$/softp�art/genl�ink?help=/md/tpKa.dgF����� �b��9�K�]�oρϓ� "Ϸ���������ߠ� ��G�Y�k�}ߏߡ�0߀�������������zQf�R�R5� ($��w���e��8�����Y  zQX���S������FH?ND[27]��!j$P��Q���Q�� � |���	����D��X�P�V���R��`  �8���ܢSB 1�XR/ \ }@�REG VE�D����who�lemod.ht}m	singl'�doub>�tripVbrowso��� �����#5�^���#dev�.s,l�Q�1�	t�}�Y� )/;/M//q/�/�/�/�/�/� tP�/? ?0?B?T?f?x?�?�?�6 @�/�?�?�?O O%O�6���/�/YOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_ �_k�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!�/ \n������ ���?"�4���j� |�3OEO+ď��я� ���+�T�O�a�s� ���������ߟ�_ ��9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}�K��ʿ ܿ� ��$�6�H�Z� U�~ϐ�_�q����Ϗ� ���� ��-�?�h�c� u߇߽߰߫������� ��@�;�M��m�g� ������������ %�7�I�[�m������ ��������&8J \n������� ���"4������ |w������ ///+/T/O/a/s/ �/�/�/w��/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?O#O 5OpO�O�O�O�O�O �O�O __6_H__�)_~_�_�Z�$UI�_TOPMENU� 1iP�QR 
d�Q�HA)*defa�ultSO<M*�level0 *>K	 �_� 5o��_3oEbtpio�[23]�(tpst[1yhGo�oWo�i/wizin?st.stm�o�&�
h58E01.�gif�o�(	me�nu5y�`*q13z)rz't4/{a��{����� �GB�%�7�I�[�m����prim=�*qpage,1422,1����я� ����+�=�O�a�s�����class,5��ß՟���4����13�H��Z�l�~������53��̯ޯ������8��O�a�s��� �����Ϳ߿���@I�P�Q�_M��]?�`a=�w��fty�m<ro�amf[0�o��}	��c[164yg�59yhae��M�#x2W-}��CzO9w {�ߋs-�?��*�<� N�`﫿������� ��m���&�8�J�\��2n��������� ��z���!3EWi ��
6����������1�0BTf�x����ainediEϯ�������config�=single&>��wintp��/ B/T/f/x/'�9Ϯ/]���gl[4�oY�H�/���!8��� 6�i�?"6�*$42h?[6��*�/G?�?3}.z>r4sx�?��8xB� <t~ۍfOxO�O�O�O �O���O�O__,_>_ �Ob_t_�_�_�_�_�_z!;$doub!%�o��13��&du�al�Y38�,4�_2oDo�_9�_n	o aVo�o�o�o__�o� 2DV%3jo=����ob8^�� ����o�"�4�F�X��+:r�Y48,2��b�ď֏�  �/�Y�k����?Y����s��v����σ�u ��N�8ߪ���?4J.�hS���w�6��u7�� ���ۯ����#��o G�Y�k�}�����0�ſ�׿�����1�"1k�}Ϗϡϳ� ����������1��� U�g�yߋߝ߯��� ����	��-�?�����6F�{������$��74ί���#�5��G��3���r��.GM?_SETUP:�������4Load� Simulat�ion�1App�ly DCS I}Ob�PTX[2˙�19MH ?VALVE ���ߙ�1/FR/C�STRT.JPG w������	A�g�CN�504JjMH��s�����"$SIN�GLE##�v381�,19 ��>26�ok}� !�y062�����/�v!��x95�Z/l/x~/�/gDOUB-�ᜃ��@ UJ/�/�??��zb `1	3��T28��?�?�_�}�treeview/4��j5i�OO %O�?�,@�?l?O�Od�O�t#2?�w93͠29 cO�O__)_ t�AO�,bO._�_�_�_�`��_�_)�GM Docs9���e�#o5o GoYoko}o�o�o��� �o�o�o'9K�o�� �O��� ���L��'�9�K� ]�o��������ɏۏ �|��#�5�G�Y�k� }������şן��� ���1�C�U�g�y�� ������ӯ���	��� -�?�Q�c�u������ ��Ͽ��ϴ_�_;� ��J�gc�k�ϛϭ� ���������u��=� O�a�s߅ߗߪ߻� ������0�B�T x��������a��� ��,�>�P���b��� ����������o� (:L^����� ���k�$6 HZl����� ��y/ /2/D/V/ h/�)Ϟ/M��/)��� �/�/	??.???Q?c? �/o?�?�?�?�?�?�? OO��NO`OrO�O�O �O�O/�O�O__&_ 8_�O\_n_�_�_�_�_ E_�_�_�_o"o4oFo �_jo|o�o�o�o�oSo �o�o0B�of x�����a� ��,�>�P��t��� ������Ώ}/�/��/ (��?-OK�]�o����� ����ɟ7�՟���#� 6�G�Y�k�}�?O��Ư د���� �k�D�V� h�z�����-�¿Կ� ��
�ϫ�@�R�d�v� �ϚϬ�;�������� �*߹�N�`�r߄ߖ� ��7���������&� 8���\�n����� E��������"�4����*defau�ltC��*level8�����������]� tpsOt[1]����y���tpio[23������u������h�z	menu7.�gif{
�13��	�5�
��
�4�u6�
��!3E Wi{����� ���///A/S/e/�w/�/"prim�=�page,74,1�/�/�/�/�/�?"�&class,13?H?Z?l?~?�??125�?�?�?�?OO#&<�?NO�`OrO�O�O�/�"18 �/�O�O�O	__&O026"_W_i_{_�_�_~��$UI_USE�RVIEW 1���R 
���_ ��_�_ym
o3oEoWoio {oo�o�o�o�o�o�o /AS�_`r ��o������ +�=�O�a�s���(��� ��͏ߏ����"� ��]�o�������H�ɟ ۟������5�G�Y� k�}�(�2����� �ү ����1�C��g�y� ������R�ӿ���	� �Ư(�:�LϾ��ϙ� �Ͻ���r�����)� ;�M���q߃ߕߧ߹� d�������\�%�7�I� [�m��������� |����!�3�E����� d�v������������ ��/ASew �������� �Oas��: ����//�9/ K/]/o/�/,�/�/�/ $/�/�/?#?5?�/Y? k?}?�?�?D?�?�?�? �?O�/�?,O>O�?bO �O�O�O�O�OvO�O	_ _-_?_�Oc_u_�_�_ �_NX