��   ~�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DRYRUN_T�   � $�'ENB 4 NUM_PORTA �ESU@$S�TATE P T�COL_��PMP�MCmGRP_M�ASKZE� OT�IONNLOG_�INFONiAV�cFLTR_EM�PTYd $PR�OD__ L �ES�TOP_DSBL�APOW_REC�OVAOPR�S�AW_� G �%$INIT	R�ESUME_TY�PEN &J_  4 $(�$FST_IDX؞P_ICI ���MIX_BG�-A
_NAM�c MODc_U�Sd�IFY_T�I� xMK�R-  $�LINc   ��_SIZc H�x� k. , �$USE_FL�4 ��&i*S�IMA�Q#QB�6'SCAN�AX�S+INS*I��_C7OUNrRO���_!_TMR_VA�g�h>� i) �'` ��R���!�+WAR�$�}H�!{#NPCH���$$CLA�SS  ����01��5��5%0V�ERS�.7  �:�6|/ 055���E����Y0�61071�5��%71�?���?d�?��_5I2j;�(O:OLO^OpO�O �O�O�O�O�O�O __�$_6_H_��FW?<N8u0 ���_��_�_����o { �2j; 4%RTNCOREV_���aL���%,o:o Ke�1(oBmo /Qo�o��'f@�o�om�o��Y�o0�� dvUx�S ��j=�9Y0�� X�r�1�tX��+01 Y0�>���,�>�P� b�t���������Ώ�� �6�1�q�1��&�8� J�\�n���������ȟ�ڟ�44�6�S!2>j9 �=� O�a�s���������ͯ ߯����/�H�Z� l�~�������ƿؿ� ��� �+�D�V�h�z� �Ϟϰ���������
� �.�9�R�d�v߈ߚ� �߾���������*� 5�G�`�r����� ��������&�8�C� \�n������������� ����"4FQ�j |������� 0BM_x� ������// ,/>/P/�