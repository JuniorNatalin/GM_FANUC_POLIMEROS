��   e�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����CELL_GRP�_T   � �$'FRAME� $MOU�NT_LOCCC�F_METHOD�  $CPY�_SRC_IDX�_PLATFRM�_OFSCtDI�M_ $BASE{ FSETC���AUX_ORDER   ��XYZ_MAP ��� �LE�NGTH�TTC?H_GP_M~ a �AUTORAIL�_}0�$$CL�ASS  �S����D��DVERSION�  ��:�8LOOR �G��DD8�?���m��Mn,  1 <DY�H8G}~}��E���82 ����D���i?/Q/@c/5/�/�/�-_ �/��/�/�+�$MNU�>A2"�d � 8iD<���?V�?V� �:�Y��MQ�L�u?��N��wQ��=�,d �80��ke?�a?�? �?�?�?�?�?�?OO %OOO9O[O�OoO�O�O �O�O�O�O�O'__#_ ]_G_Y_{_}_�_�_�_ �_�_o�_oGo1oSo }ogo�o�o�o�o�o�o��o	U?7N_UM  ��>a� �p���2T�OOL?#8^�����%>�n��:���?�����Q���nn�:����p�����£�C���Mv\gŽ��o�?!�<����?�=���� �Y��?\TB�����}U�D�D9Mva^-�{�Î>�<��j?���kr��<y���?ae�C�l':�D�Kx^����qfqeu�p��|�B��\)�y��DS������#�!+�Oq�����'����e�����>���C�&A��-�?�9�dż��>�U<`���?�;�����6T���?ak�����s�{q�C�/�S�e�������O�@�{�G������B����~ffB��� ����ﯡ���%��1� [�E�g���{���ǿ��@����ϭ�v�s[�y 