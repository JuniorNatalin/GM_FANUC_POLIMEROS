��   ��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����PMC_CFG_�T   � �$'NUM_MS�K  $EX�E_TYPECM�EM_OPTPN�_CNFCIF_�CY:gSCN_�TIME E R?ESET_P�D�o LJ �HECK�_DSBLC $�DRA> ARGI=NCSTORJ2 �&DEV. d� 	7OC'HA�R�ADD�SI�ZORACBSLmO[ODKIOKOCCPYC&l >/  L ��ph99IDX��d&L. � �
�EQPLHR�AT�TRKBU�F| ��UN_�STATUS�C�U��MAX(I�� �SNP�_PA�  �� � ANNE��� OW CTIO�N_�PU� �  $BAU}D�NOISYm�N�T1�#2�#3n�$_PR�T4P�' DATA�CQ�UEUE� PTH�[$MM_��%&!R�ETRIESCAUTO!R[���BG � �ISP_INFd�' C�LIMI� B5AD_H C3H��#d6�# d6�#d6�#W1� �#�4�#�4�#�4�"�� ��$$CLASS  ����1������0VERySg �8�07�:�iFG0 �5���
@+A�2��� ��d��3CC��  2G'@d $)DxO��uO�O�O �O�O�O�O__:_)_ ^_M_�_q_�_�_�_�_ �_�_oo6o%oZoIo ~omo�o�o�o�o�o�o �o2!VEzi ������
�� .��R�A�v�e����� �����я���*�� N�=�r�a��������� ޟ͟��&��J�9� n�]���������گɯ ���"��F�5�j�Y� ��}�����ֿſ��� ��B�1�f�Uϊ�y� �ϝ����������	� >�-�b�Q߆�uߪߙ� �߽�������:�)� ^�M��q������ ������6�%�Z�I� ~�m������������� ��2!VEzi ������
� .RAve�� ����/�*//�N/=/R,CIF 2]aKP )DX5D��)G�&Ȫ'�%Y��(�(�!�%� �&D�6C�9@  '^/X/"?K?F?X?j? �?�?�?�?�?�?�?�? #OO0OBOkOfOxO�O �O�O�O�O�O�O__ C_>_P_b_�_�_�_�_ �_�_�_�_oo(o:o co^opo�o�o�o�o�o �o�o ;6HZ �~������ �� �2�[�V�h�z� ����������
� 3�.�@�R�{�v������ß��П���#TY�PE 2�+ �(�#	0d�ʙ���!�����h���	0��ɯ	0ฯ���~#SNP�_PARAM ��+���1' C�q���!ۤ�"��1	0UD��)R�