��   L�A��*SYST�EM*��V8.3�382 5/9�/2018 A� 
  ����CELLSET_�T   w�$GI_STYS�EL_P �7T  7I�SO:iRibDiTRA�R��I_INI; ����bU9ART�aRSRPNS1TQ234U5678Q�
TROBQACKSNO�� )�7�E�S��a�o�z2� 3 4 5 6� 7 8awn&GINm'D�&��)% ��)4%��)P%��)fl%SN�{(OU���!7� OPTNA �73�73.:B<;}Ta6.:C<;CK;CaI_DECSNAp�3R�3�TRY1���4��4�PTH�CN�8D�D�INCYC@HG�KD~�TASKOK� {D�{D�7:�E�U: �Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T�8�T�@REQ�d��drG�:Mf�GJO?_HFAUL�Xd8�dvgALE� �g�c�g�cvgE� �H�dvgNDBR�H�dg�RGAB�Xtb �Z �CLMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVERSION�ix  ��:�$'61�r���p��q�t+ �UP0 �x�Style Se�lect 	  ���q�uReq.� /Echo��N�yAck�����InitiaQt�p�r�s��#��@�O�a�p���	���  ����*������)���������q���O�ption bigt A��p ��B���C���Decis�c�od;��w�pTry�out mL���
�Path s�egJ�ntin.z��8,� cyc:���\�ask O�K!�Manual opt.r�pA"��ΜB"�#�Μ�C"�?�Δdecs�n ِ��pRob�ot inter�lo�"�<� i�sol3�"�̕CҚ�i/�"�x�ment��x�ِ���"���^�statu�s�
	MH ?Fault:��'�{�Aler��ǁ'���p@r 1�z L��[�m�+��; LE_COMN�T ?�y� � ����������ۿ� ���"�4�F�X�j�|� �Ϡϲ����������@�0�ƿ@�>���s�25 ��Too�l Change<��*�
Cap���_Auto ��r{��y��Repai������2�r3���
��4��Re�served��'�BY�cW諸80�373 ��� '�tm������hᦈ������z!��i��bI��G�H���Gw��;(
�������֚�<��(���m�� C%(n��N9"�&mKu(�M��� �R�(Ҷ��� mZ)��)� $Qae)6�=y )�mi�)h�H�� .�p/)�n.Zz/�A/�xU/)�-/��i/�/��/)m�}/޹/�/���/*0�/�	?1>H��0b�?\U� %�? mR�? ��? *�?� :�? G�? Ơ�?�?�?O���IO ud]O �?  [�O4GO�p4�O h�O�O4�O�]�O i_Sߢ�p�9_7_�p�a_ ��Y?+�ZD�T Tes����t�eBreakΫ�eck��nc�l�_+��^
udv�_ �ncesom,d
v�  �/�T fQo,V=oimoyo ��_de�o�,��ou/  �X�n.p�o,��oUX?\l�A~��A,�/7
EBi W?�  -}�Ġǈ���pP��Ġ� 1�/��p�/.����V�"�q�m���Ġ�яϏ�p潏��Ġ�/��!��G�ĠPF�!J@]���Ġ����!|��D�Ġ��� ���D7�Ġ�a�_� �M�䇯�������  /���ׯ0 � �/D���0��֯Z�v=�35y����***��/���]�ɿ��ǿ��ݿ4? �Ϙ�m00?
�� ;
<o 0>}�gϺ0!U~$NU��0h�oN�1&U~�xh� 0��REY��+U~EG/ 0Ժm�s�� 1U~tm l? 1d�
iL� �8.2!�1E8�d o����h�o� 1j]�o�0� �f�o 1���*]F��G�o@��!/ߣ K�u���D'� � ,�$STY�LE_COUNT�" ��������ENAB  �������� 0������� ���	����DV k����� �,>P�q ��������� //(/:/L/^/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�?x�?�=��MENU������6NAME ;?%��(%f�B�_��IO]UY%	P�RT03_R02D0O7I$EVO^O5qOD3MkB6�O�Om@7�O �O�O�O1_j_U_�_�K#11_�O�P2�_�_ �PpO"_�_5o oYoDo }o�]_�_�Q8�o�ob�P9�b�o�L20�o ouo�oAJm0Bdo��%d�h2Odv� ���-�?�Q���u����YxMOV_REPR���Ё�o�Ё)3����4.����@�d��9h������r��˟>�kA3p�o����� 
�C�ޖ4�_�o\��_"� [� o2�4��Я	���p�O��������J���.���ښ5:���@����!���E��:�Ds�!�9bϛ�	�L��D��!�>����	�~��D�!�D�;�	�*�Dc�!�IRߋ�	��z���!�O����  2���!�T��+���F�S�!�ZB�{���xj��!�`�����������!�e����Б�
�C�&�k2�k� G 3Z���&�q��D��~�@����&�v��D~�r��3&�|"D[~�J�&ЂrD�~�֚�&Ї��  4�#&��K::s&��b�l��&������/&�/:/�*/c/&�q��/�p5z/�/&Щ��/�/� 4�/?&Я��/+?� f?S?&д�B?{?� ���?&й�%�2101_TCɿ�w�52�?�?�03�?�?�04O&O�05<ONO�06dOvO�07�O�O�08�O�O�0y9�O�OE110_�޿�2-T1_  6� J_�_F_�_jT��_�_��_�7(�_#o&Ё�oKo`i�ro%��bo�o`��o�o&���o�o`��o&��Y 4g�ob%��R��&�gz� � ��%repair��\�328_Z#DT��W�t9��_� ̈B�{�6ϟ��� Q�ʏ�qY쏇���� �
�C�&��	�j�����no����&�<���~�� ���(�:�L���p�����ͯ�a��P#:H�#��?�K�"�z:�s��Eb���"����ÿ�J�����ڿ����:�P;*�c����M��Bzϳ��ao��M�t�����_��+�N��@�S��	�z�M��j����j����  <
�����p����ЈџB��u2�k���n�Z���{����Р�����栀���������3�栆"�[�  =J���栱o��m�6����树����n�h��#栗Kn��:s栝b�n�̊�栢��n���栨; G >0*c栮RD�Nbz�栳�D�N��/根�+/N�/S/�z/M�j/�/���/P#?*�/�/���/?"� \
?C?��2?k?"� �Z?�?�Ղ?�?"� ��?�?���?O"� ��?3O��"O[O  @$JO�O�9o�OmAV�O�O栉o�O�mAi�"_�QJ_mA�:_s_��b_�_���_�R��_�_  � �_o�_5o!d(oao$o�oqd�xo�oto�o�f�o�o'. 6HZl������tLE���r
�C�ΐ�2�k�.���z� ��ި�o⏥���� �'�9�K����p����q���ӟn����r�.�=�#� yq�K�  �:��s� FIb��� �O��¯  MEyN��� )�گ �����:�L`D	�b�2��`R��� !蟱��L`����ڿ  &y�