��   X�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����CIPS_CFG�_T   0 �$INTERF�ACE  $�DUMMY1B2rB3B&SET/� @ $MO�DA8 _SIZ�}OUT�DAT�E_FIX~CS�I_VRC  �  ��$$�CLASS  O������O���O� VERSIO�N�  �:�$'1 �O� �m r �
��� � /� -@