��   ~�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DRYRUN_T�   � $�'ENB 4 NUM_PORTA �ESU@$S�TATE P T�COL_��PMP�MCmGRP_M�ASKZE� OT�IONNLOG_�INFONiAV�cFLTR_EM�PTYd $PR�OD__ L �ES�TOP_DSBL�APOW_REC�OVAOPR�S�AW_� G �%$INIT	R�ESUME_TY�PEN&J_ � 4 $(F?ST_IDX�P�_ICI�T��MIX_BG-<A
_NAMc gMODc_USd~�IFY_TI�w �xMKR-�  $LI�Nc   �_SIZc�x� k�. , $USE_FL4 �p�&i*SIMA��Q#QB6'SC�AN�AXS+IN�S*I��_COUN�rRO��_!_TMR_VA�g�h>�i) �'�` ��R��!�+W[AR�$}H�!�{#NPCH���$$CLASS ? ���01���5��5%0VERS��.7  ��:�6/ 05�5�������Y0�61071�5���%71�?���?�?���_5I2j;  �?9OKO]OoO�O�O�O �O�O�O�O�O_#_5_0G_��FW?N8u0� ���Z��6�[�\ @�Z	��L�o { 2j; 4%V_o����1�1�_9o diqroao��>
<Po�o��:CO�o�o���ent�o�o��T��o1C"g���̀Ty�S��j=�9Y0`�� �r�1�tX��01Y0�>���,� >�P�b�t��������� Ώ{�5�1�q�1�� &�8�J�\�n������� ��ȟڟ�44�6�S!�2j9  �=�O�a�s������� ��ͯ߯����\/� H�Z�l�~�������ƿ ؿ���� �+�D�V� h�zόϞϰ������� ��
��.�9�R�d�v� �ߚ߬߾�������� �*�5�G�`�r��� �����������&� 8�C�\�n��������� ��������"4F Q�j|����� ��0BM_ x������� //,/>/P/�