��   �=�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����EIP_CFG_�T   � �$VENDOR � $DEVT�YPE>PRDC�ODIREVIS�ION>FAST�_UDP 5 K�EEP_IO_A�nSCNpOPT�` Sp $LOAgDED� �CC� �IG�ED_MO�D�NET�EX�PLCIT_MS��$HIGH_�SPEE�$E�N8021pDS+CP� Hp �� �SPARE���&ONN. |� $HOS� �!B SC9ENA�BL$STA�TN _SZ�S�^TOAPI�OETrIgA�R]�V�BW&Mo� &SC.�  7�CXQ�[XX_���CX_��[ kRs�)%'FLA�MU�L�TR�� C_�O�["TOD&IC$i �AS�Z 'sEC{#�#TIMV�CN� Z�&PAT�  @$IDA_FORMA���!�&� �"9"FIG�^�"2�+�!�$ANALOGI� o  4OU� f8FM�$Q�(���$$CLA�SS  ����e1��.��.Z0V�ER_c7  �:�$'�0 �8. d����0�0> �?�1�1���7/ ��4(� 2�;@ p!�124.11.�240.31�����1  [2�5;��P!Ce�ll ctionPABO�6�12_D<gD��:!l1�O��!Conne:BbA�O�OKOyO�O�O3_1_C_�Og_
_<@4q_�_�_V_�_z_<@5�_o#o�_Go�_<@6Qo�o�o6o�oZo<@7�o�o�o'�o<@81as�:<@9������<@A�A�S��w��<@B����Ïf�珊�<@C�!�3�֏W���<@Da�����F�ǟj�<@Eџ����7�ڟ<@FA�q���&���J�<@G���������<@H!�Q�c����*�<@I����ӿv�����<@J�1�C��g�
�<@Kqϡϳ�V���z�<@L���#���G���<@MQ߁ߓ� 6߷�Z�<@0���ߖ���)���nO1�a�s���:�<@P�����������<@Q�A�S���w��<@R������ f�����<@a0#����Y��nTa��F�j<@U���192.16�8.1C?�@Ou�tputVlv#<QN�8�;���L�W����/��A3_K/]/ 2�_~
#
MH InX ^o}�,�_�-�O /?�/�/6oo�-:/�? B?��?(/�oOO / AO�?6!O{O�O0O�O TOfA��O�O�O!_�Of@401_\_n__�_ 5_GP�/�_�_�_o�_ FQ?;oMo�_qooFQ �?�o�o`o�o�oFQ�/ -�oQ�oFQ�/� �@�dFQl?�� �1��FQ�?k�}� � ��D�FQjOۏ폐�� ��FQ�OK�]� ���$�f@5J_��͟p�񟔟 ���_+�=���a���� *o����P�ѯt����o���p/25
��D�KL ChangSerQ�r̠+� ɯ����z�����!� Ŀ���[�m�ϑ�4� ��Z����π�ߤϦ� ʏ;�M���q�ߦ�:�@�߽�`��߄�f@6�� �-���Q������� ��@���d�ኯ��� ��1������k�}� ����D��L���������$EIP_SC �2����. @������ K����[@ ]�����}r���,>P bt������ �//(/:/L/^/���:�/t/�/�/�/@ Rdv'?9?K?�o? ��?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�O�O�/_ _C_U_g_y_�/�/? �_�_�_X?�_|?-o?o Qocouo�o�o�o�o�o �o�o);M_ q��,_>_��� ���_�_�_�_m�� ��ooǏُ���� !�3�E�W�i�{����� ��ß՟�����/� A��e�T������� � 2�D�V���+���O� s���������Ϳ߿ ���'�9�K�]�o� �ϓϥϷ�����r��� ��#�5�G�Y�̯ޯ� �߳���8���\��� 1�C�U�g�y���� ��������	��-�?� Q�c�u��߈����� ����f�xߊߜ�M_ q���ߧ���� %7I[m �������/ !/��E/4/i/{/�/  $6�/�/?~/? �S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�OR/�O �O__'_9_�/�/�/ �_�_�_?~_<?�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CU�O�Ohz� ��F_X_j_|_-�?� Q��_�_��������Ϗ ����)�;�M�_� q���������˟ݟ� ��%��I�[�m�� ���ǯٯ�^�� ��3�E�W�i�{����� ��ÿտ�����/� A�S�e�wωϛ�2��� �������ߌ����� a�s߅���^������ ����'�9�K�]�o� ������������� �#�5�����H�Z��� ����&�8�J�\� 1�߶�gy��� ����	-? Qcu����� �x�/�)/;/M/�� �������/�/�/>�/ b?%?7?I?[?m?? �?�?�?�?�?�?�?O !O3OEOWOiO{O/�O �O�O�O�O�Ol/~/�/ A_S_e_�/>_�/�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o�O�O(:o ��__*_<_�� ��_�_G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��X�ԟ	��-�� ����������ϯ B����)�;�M�_� q���������˿ݿ� ��%�7�I�[��� nϣϵ�����L�^�p� !�3�E߸��ܯ�ߟ� ������������/� A�S�e�w����� ������Ϟ���O� a�s�����
������ ��d�v�'9K]o �������� #5GYk}� �8�����/�� ������g/y/�/���/ "�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;O�_O NO�O�O�O�O,/>/P/ __%_�/�O�/m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�olO~O�o�o/ AS�O�O�O�O�� �D_V_��+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ������ɟ۟�` r��G�Y�k���� ���ůׯ����� 1�C�U�g�y������� ��ӿ���	�ϲ�?� .�c�uχϙ���0� �����x��Ϝ�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ����L�^������ !�3��ϸ����ύ��� ��$�6�����/ ASew���� ���+=O a��t���@� R�d�v�'/9/K/��o/ ���/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?�?�?�?�?�O OCOUOgOyO��/ �O�O�OX/�O|/-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o,O>O�o�o�o �O�O�O�Om �__����� !�3�E�W�i�{����� ��ÏՏ�����/� A��oe�T�������  2DV��+��O� �s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿr��� �#�5�G�Y�̟ޟ� �ϳ���8���\��� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u��ψ��������fψ��	��4��� $i,�,d��b�t����Ϫ��� ������(:L ^p������ � $��H7l ~��u�'����� /����)/V/h/z/�/ �/�/�/�/�/�/
?? .?@?R?d?v?�?�?�? �?U�?�?OO*O� ����O�O�O/�O ?/�O__&_8_J_\_ n_�_�_�_�_�_�_�_ �_o"o4oFoXo�?|o ko�o�o�o�o	�[O�j>:�j,h,gBT�C�o�O��� �����!�3�E� W�i�{�������ÏՏH����l�|O
� � R�d�v��on-�|� ����Oy*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ����;�ȿ�o���� ����7Ϲ�˟|ώ�� �����������0� B�T�f�xߊߜ߮��� ��������,�>�տ b�Q�����OOA� sO��(���L���p� ��������������  $6HZl~� ����o���  2DV������\� ��G�Y�
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�? cu��JO\OnO� ��O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo�? Bo1ofoxo�o�?O!O 3O�o�o{O,�OP bt������ ���(�:�L�^�p� ��������Oo܏ˏ � �$�6��o�o�o<��� ����'9���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�����w�����п C�U�g�y�*�<�N��� ӟiϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶��������ߕ� "��F�X�j�ݿ�� �������[���0� B�T�f�x��������� ������,>P bt��/��� �����p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?�h?W?�?�?�? #5GY
OO.O� �IOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_u? o�_&o8oJo�?�?�? �?�o�o�o;O�o_O "4FXj|�� �������0� B�T�f�x�o������ ҏ���io{o�o��P� b�t��o�o����Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$���H�7�l�~��� ��'�9����ρ� ��)�V�h�zόϞϰ� ��������
��.�@� R�d�v߈ߚ߬߾�U� ������*���� ӿ�������?��� ��&�8�J�\�n��� �������������� "4FX��|k� ���I�[�m��0 BT������� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/?�(??L?^?p? ���?�?�?a s	O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_5? �_�_�_�_
o}?�?�? �?dovo�o�?�oO�o �o�o*<N` r������� ��&�8��_\�K��� ������)o;oMo��� "�4��o�oj�|����� ��ğ֟�����0� B�T�f�x��������� ү�{����,�>��Pf�̇�x�	��4�� $�,d�,e\�¿ԿG�� H�d��'�9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}�������������� ɏ{����P�b�t�G� ������������� (�:�L�^�p������� �������� $�� H7l~���'� 9������)V hz������ �
//./@/R/d/v/ �/�/�/�/U�/�/? ?*?�����?�? �?�??�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_�/|_k_�_�_�_�_ I?[?m?�_0oBoTo�? �?�o�o�o�o�o�o�o ,>Pbt� ��������_ (��L�^�p��_�_o oʏ܏�aoso	�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�����5�¯��� ��
�}�������d�v� �������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�ϯ\�K߀ߒߤ߶� )�;�M����"�4刺 ��j�|�������� ������0�B�T�f� x�������������{� ��,>P������ �ߪ��A�S�� (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/ �/�/]o��D?V? h?��?��?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _�/<_+_`_r_�_�_ 	??-?�_�_oo�? �?Jo\ono�o�o�o�o �o�o�o�o"4F Xj|����[_ ����