��   ,��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DCSS_IOC�_T   P �$OPERAT�ION  $�L_TYPBID�XBR1H[ S2�]2R �$$C�LASS  �������P��P�� VERS?��  �:��$' 2 ��P @ �����  
�*����	��� ���������� ����V ��f"Nj>�������� ~����F��b��� :!�
!J�F�� ���/����@��������/ 1��/  �S(��?  ��^)������
/  �&/ s �B/  �N�  �z/ ���  �V���sO �֏O  ��O !��1�"�61�#��R1�$�n1�%���1�&��1�'���1�(��1�)���1����A�+��2A�,���-��jA�.��A�/���A�0��A�1�C"? � D>?  �3C�4Cv?  95�4�o  6�4�o�  7�  8 �.}u��������_C_CCL �?��  �	All par�am��
Bas�e�Pos.�/Speed c�heck(�Saf�e I/O co_nnect�}R���pConfig�ChngRese�tTotal�0����1�0�-S�p��, Onn�wS�Ii�@�pNoGenStopN���ypas�No�Es��0Fen�ce Statu�$��1��rved���D�V�h�z�E�xtS��oDisbl4�}�������ŏO��n����'�9�K�����CPCZo3ne�av�ne�a��3ne�a��ne�a��3ne
q֯ne&q�3neBq�ne^q�ne9�~�~aO�e1��T���T���T� ҦT��T��T��T�2�T�J�T�2c���{� ����������ÿ��ۿ ��󿝣ϝ�#ϝ�;����Sϵ�kϵ���Jo?intChk[݃ՠs߅ӛ̓ճ�~�artSpd���ޢ��~���S�e5��=�2�N�J�N�6C�}슧~����~뺧~�ҧ�|SO<��pNo �V�}
��s OFF
��Teach;� OAutoL�M�T���e��M�Enba�bleDevic�e��H�ty�w�orkActiv�蓩� dis�� �switP�-���Ma��͔���唏��� 0�5������U�d�^��GYk^Ճ�4��2 ����ͣ�������-�5E�M [�4�s�s�s� s�sss4 sLsds2}e� n/~Æ/�Þ/�ö/�� �/���/���/�?&� .?>�F?V�^?n�v<�ր�?�Ӧ?�Ӿ?��v; ��4���=6��H +O$C<�N�gOr����O��������C_N揅`����;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ ���������ZSIh���IO� Interlock3�"��}����� ��ŏ�����6�1� C�U�~�y�����Ɵ�� ӟ��	��-�V�Q� c�u����������� ��.�)�;�M�v�q� ��������˿ݿ�� �%�N�I�[�mϖϑ� �ϵ���������&�!� 3�E�n�i�{ߍ߶߱� ����������F�:��P%_�24Vo�utaftMCC���NonMtnBreaker��SFDI�M��]��5���6���cM ��{M?�G�3�E�W�n� {��������������� /FSew� ������ +=Ofs��� ����//'/>/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?^? k?}?�?�?�?�?�?�?��?OO6OCON�`�OHd�8P��O�M�O�M �E��C���C���C�� �C��C&�A�Q_c_�_ �_�_�_�_�_�_�_o o)o;odo_oqo�o�o �o�o�o�o�o< 7I[���� �����!�3�\� W�i�{�������Ï� ����4�/�A�S�|� w�����ğ��џ�� ��+�T�O�a�lO_��Sc��BVOFF~n�FENCE��?EXEMGկ�����NTED��OP��AUTO�T�O[��O�|����CSBP蔿���Ov�No� General� Stopǧen�ce ԭ߰E�xtern�E-��߰Serv�o Discon�nect|�C_D���_`�S�y� 