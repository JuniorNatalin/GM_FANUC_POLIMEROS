��   �A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����FSAC_LST�_T   8 �$CLNT_N�AME !$�IP_ADDRE�SSB $ACC�N _LVL  �$APPP  � ��$8 AO  ����z�����o VERSI�ONw � �:�$'DCEF\ w { �� ����ENABLEw �����LIST 1 �  @!�$�����
[ .@�d���� �/�3//W/*/</ �/`/�/�/�/�/�/�/ �/??S?&?8?J?�? n?�?�?�?�?�?O�? �?OO"OsOFO�OjO|O �O�O�O�O_�O�O7_ _\_B_�_f_x_�_�_ �_�W