��   �i�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DCSS_CPC�_T   � �$COMMEN�T $EN�ABLE 6 M�ODJGRP_N�UMKL\  $UFRM\~] _VTX 6 ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�?  &S. Ǆ 8J\TC��u
SPD_LI`_���SOL��&Y0  � �1CHG_SIZ�$APGE.SDIS��GB�C����J
p 	�J�� &��"�))$'2_SyE�� XPANI�N��STA�T/ D $�FP_BASE �$_ K�$!Y �&_V�.H�#�  �&J- q�ZAXS\7UPRJLW7S<e� x��$� | 
�/�/�/�D&?8?z�&EL�EM/ T ��2�"NOG�0�3�UTOOi�2HA�D�� $DAT=A" 0&e�0  @@p:�0 _2 
&Pp%' � p!U*n   �FS�Cz�B�� �B(�F�D(�R|UC�DROBOT�H��CqBo�E�F$OCUR_2R &�SETU�	 l|� �P_MGN�INP_ASS� 0"@�� �3�8B7gP@@U�^V�Sp!��&T1�
`B|8�8�TM 0 6P�+ Ke�1VRFY�8
dD5F1�� ��W��1k$R��&TPH/ ({ �CA�CAt�CA3�BOX/ 8�0����У�b'oEcd�TUI}R�0  ,{ �FR`ER�02 {$�` �a�_S�b��fZN>/ 0 {9F02� -a0rZ_0��_0�u0  @�Q�Yv	�o:n ���$$CLLP  O����q��Q���Q�pVERSIO�N�x  ��:�$' 2� �xQ   �Press��8���p� �p�q����#PE��� ņ`�1�D?/  E��M���B�����
�� ��
Tool C�art ��)�;�Z�� EC�U��;�g C��z��Ȉ�2 ��� �qJ���ˏ�9���]�����R� ����g���������9� _�q�������L�:��̯����Fen�ch By Pl?atformU�g�~y�g@ Ň�����
����s��)H����0�e5���࡯O�a����W� �z%���*�!�״onveyor�@��y���������\����� ���φ�'ߪ� ��/���mߓߥ���� 8�J߀�n� �5�G�� k�����"������� X��|���U���y� ������0�B���f� -��Q<����� ��>�t� ;�_q�� (�L//%/�I/ ��/��/�/�/6/ �/Z/l/�/�/1?W?i? �/�?�/?D?2?�?�? Oz?/O�?�?�?wOfO �O�OO�O@OROdO_ �O=_O_�Os_�O�O_ �_*_�_�_`_o o�_ �_]o�_�o�oo�o�o 8oJo�ono#5�o�o k�o�o���� X�|�C��g�y� ������0���T��� �-���Q���ҏ��� ����ϟ>��b�t��� ;�*�_�q������� (�ݯL�����7��� ��ʯ����$�ٿ ĿZ�l�!ϐ�E��ƽ��$DCSS_C?SC 2�����Q  Dֿ��f�˘��ϼ� ��#���5��k�:ߏ� ^߳߂��ߦ������� 1�C��$�y�H��l� ������	���-��� Q� �2���V���z��� ��������;
_�.@��v	�z�G�RP 2�� 	���	<�!E 0iT�x��� ��/�///S/>/ w/b/�/�/�/�/�/�/ �/??=?(?a?L?�? �?�?t?�?�?�?O�? 'OOKO6OoO�O�O^O �O�O�O�O�O_�O5_  _Y_k_}_H_�_�_�_ �_�_�_�_o
oCoUo go2o�ovo�o�o�o�o �o	�o-?Qu `����������_GSTAT� 2���,8��?w����TT?>~����Vs<��  ���ewb���a�ҿ[�E�ü�YD�s�����8V�k��g�.��,���4���Z��j���D4  ��"�����V�����M6�,n?�w6�׀7^I�(΁��Cۥ��D��|ƅ��]X 5W��?�7bo������9��W�J�7C����n{D�����ϵT���g���&��gxj�=�a�Eሼ�?�'D��pƅZ��c%b�7f(ؾ��5��=�s�6#?�Z�b�X�j�|� ����������(�:� �^�p���	ɒ��n� ��ͯ��ɯ����� #�5�W�Y�k�����ņ v��B��&�8��\� nψ�¿�Ϟ����ϸ� ������:�$�F�p� Z�lߦߐ�N������߀�0��T�f�D箐����J�>~�ﶜ�x�����'��5I��ΐ��~��� �D�{rq����l���+�����Ᲊ��Ex�a5�X�cր3ڀ36���5����Cۤ����Db��z�� �4����	6���Q��Q�=��m2�#C� ��׻Xm2��*���s�:�J�D�R�ﶋ�ྒ������y�D���K~�>���6�� ����㈾�������� ���J�.Rd B���Ϻ����� ��0,fP b�����z/ &/xJ/\/:/�/�/� ��/��/�/�/�/? ?$?F?p?Z?|?�?�? �?�?/OOp/BOTO 2OdO�OhO������� ��������(�:�L� ^�p����������_�O �O �OLo�O<o�o�o ro�o�o�/�?�o�?  *6`Jl�� �������oD� V�4�z���j����o �����"��.�X� B�T���x��������� ����<�N���r��� b������O
oo�O�O �O_"_4_F_X_j_|_ �_�_�_�_�_�_�_� ��0oj�|ϖ��ϲϐ� ����Ώ���$���0� Z�D�fߐ�zߜ��߰� �������2����t� ��d��������� F��"�(�R�<�^��� r��������������� *��l~\�� ���ԯ:�L�
�� .�@�R�d�v������� ��п����� &`Ϛ/�/��/�/�/ ??��(B?L>?`? b?t?�?�?�?�?�?�? O,OO8ObOT�O�O �/�O�O�O�O_*?<? vOL_ROX_�_l_�_�_ �_�_�_�_�_$oo0o ZoDo"_�o�O�o�o�o �oX/j/|/:L ^p������ � /J/$/6/H/2D V�oʏ܏�� ���� 6�H�._hor�|o~��� ����ޟȟڟ����� 2�\�F�h����o¯ԯ &���
��.�@�Z��� j���f���������� ҿ����*�T�>�`� �ϰ����������� �8�߈�����j| �������� �0�z�T�f�l�b�t� ��(������0�B� � f�x�^��Ϣ�tϮ��� ������D.@ zdv��X�� �(:^p��� ������/� /$/&/8/Z/�/n/�/ �/��/�/N ?2?? V?h?R߸���ߚ߬� ����������*�<� N�`�r���O�?�? ��x?*_|?:_`_>_P_ �_�_��/�_�/�_o �_o>o(oJoto^o�o �o�o�o�o�o�_"4 XjH���_�o ��o� ���6� � B�l�V�h��������� ��,�
�P�b�@�������u�$DCS�S_JPC 2��uQ (G D������ ��0ԟ)���
�_�.� @�R���v�����ﯾ� ��7���m��N� `�����������̿!� �E��i�8ύ�\�n� �ϒϤ϶������� S�"�w�Fߛ�j�|��� �߲���������a� 0��T��x������ ����'�����o�>� }�b������������� ��5G(}L^ p�����1  U$6�Zl~ ����/�?// c/2/D/�/�/z/�/�/ �/�/�/)?�/M??q? @?�?d?�?�?�?�?�?��?�?7OOEO���S
��Ý@0O�OTO&O �O�O�O�O!_�O_W_ *_<_N_�_r_�_�_�_ �_�_o�_oSoeo8o Jo�ono�o�o�o�o�o �o'a4F� j|������ ��]�0�B�����x� ��ۏ����ҏ#���� Y�,�g�P���t���ן ����Ο���U�(� :�L���p���ӯ寸� ʯ��?��c�6�H� ��l�����ῴ�ƿ� ����_�2�Dϕ�h� zό��ϰ����%��� 
�[�.��Rߣ�v߈� �߬�����!����W��*�<�pHMODEL� 2�Kx�Tool Ch�anger��
 �<v�cz���CݯK� N�ĉ/� C�L�D������I���5���0� B�T�f����������� ������g>P �t�����D�����p�Y k}�����$/ �//1/C/U/�/y/ �/�/�/�/�/�/�/	? V?-???�?'9g?y? �?a?�?�?.OOOdO ;OMO�OqO�O�O�O�O �O_�O_N_%_7_I_ �_m__�_�_�_o�? �?�?�_o�_EoWo�o {o�o�o�o�o�o�o�o X/A�ew� ������B�� +�=�o��7oe�w�M� ��͏���P�'�9� K�]�o���Ο����� ۟����#�5���Y� k�������������� ۯ�Z�1�C���g�y� ƿ����������D� �-�z�Q�c�u��ϙ� ��������.���)� ����#�Q�c��ߧ߹� �������%�7�� [�m��������� ��8��!�n�E�W�i� {�����u��������� F/|Sew� �����0 +=Oa���� ����//��t/ =/O/�/�/�/�/�/ �/�/:??#?p?G?Y? �?}?�?�?�?�?�?$O �?OZO1OCOUO�OyO �Oa/s/�/�O�O2_�O _-_?_Q_c_�_�_�_ �_�_�_�_�_oodo ;oMo�oqo�o�o�o�o �o�oN�O�O) ;�#����� &���\�3�E�W�i� {���ڏ��Ï���� ��/�A���e�w�ğ _q��������� f�=�O���s���ү�� ��ͯ���P�'�9� ��]�o���ο����� ۿ�:�՟���'�9� �}Ϗ��ϳ������ ����1�Cߐ�g�y� �ߝ߯���������D��-�z�Q�c�u�K� � TI TOOL� CHANGER dϒ��������� 0�B���f�x������� ��������C,y Pbt����� �-P�b�� p����/�� ;//$/6/H/Z/l/�/ �/�/�/�/�/�/�/?  ?m?D?V?�?>P~? �?�?x?�?�?EOO.O {OROdO�O�O�O�O�O �O�O/___7_<_N_ `_�_�_�_�_�_�_�_��3�$DCSS_�PSTAT ����Aa�Q    � �0Zo`b  bn(to�o�ol�odo �k  `�B`�ar`o$�9�cAeN�`Cu~2dSETUP 	AiGB�d�3Va �t�-iT1SC 2
4�z�`�1Cz�3�����uCP R�|��0D�?X�j� �?��������֏��� ɏ�0�B��f�x�G� ������������ן ,�>�P��t�����g���ί�3��7F��� ��9�K�]�,������� t�ɿۿ���#�� �Y�k�:Ϗϡϳς� ���������1�C�� g�y��?����H��� ��	���-�?�Q� �u� ���h������� ���;�M�_�.����� ��v���������% �ߞ�[m����� �����!3E i{J\��� ��/�//A/S/"/ w/�/�/j/�/�/8J ??�/=?O?a?0?�? �?�?x?�?�?�?�?O 'O�?O]OoO>O�O�O �O�O�O�O�O�O#_5_ G__k_}_�/�/�_�_ L_�_�_o�_1oCoUo $oyo�o�olo�o�o�o �o	�o?Qc2 ���z���� �)��_�__�q���� ������ݏ��Џ%� 7�I��m��N�`��� ǟ������ޟ3�E� W�&�{�����n�ïկ <�N�����A�S�e� 4�������|�ѿ��� Ŀ�+����a�s�B� �ϩϻϊ�������π'�9�K��o߁�P���$DCSS_TC�PMAP  ������Q_ @ \�\Х\�\���\��\�\�\�	�� � \�\�\��\�\�\�\��\�\�\�\�J\�\�\�\�\�U\�\�\�\�U\� \�!\�"\�U#\�$\�%\�&\�U'\�(\�)\�*\�U+\�,\�-\�.\�U/\�0\�1\�2\�U3\�4\�5\�6\�U7\�8\�9\�:\�U;\�<\�=\�>\��?\�@��UIROw 2�������� ��$�6�H� Z�l�~�����������@���� 2[��� [������� ��!3EWi {���<�`� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?�a?��?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O�T?�O��UIZN �2��	 ��� ��._@_R_W�)_~_�_ �_e_�_�_�_�_o o 2o�_VohozoIo�o�o �o�o�o�o
�o.@ Rd'��i{� ����*�<��`� r���G�����̏���� ��׏8�J�\�+��� ������y�ڟ쟻���"�4��O��UFRM� R�����8 _ߌ���]�¯ԯ���� 
��.�@��d�v�Q� ������п⿽��� �)�N�`�w��ϖ�5� ���ϧ������&�8� �\�n�Iߒߤ�ߵ� �������"���F�X� o�|��-������� �����0��A�f�x� S������������� ��>Pg�t�% ������( :^pK��� ��� //�6/H/ _V/~/�/k/�/�/�/ �/�/�/ ?2??V?h? C?�?�?y?�?�?�?�? 
O�?.O@OW/i/vO�O 'O�O�O�O�O�O�O_ *__N_`_;_�_�_q_ �_�_�_�_oo�_8o JoaOno�oo�o�o�o �o�o�o"�oFX 3i��{��� ���0�B�Yof�x� �������ҏ䏿��� �,��P�b�=����� s���Ο����ߟ(� :��