��   O�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DMR_GRP_�T  � �$MA��R_DO�NE  $O�T_MINUS �  	GPL�N8COUNP �T REF>wPO�OtlTpBC�KLSH_SIG�oSEACHMS9T>pSPC�
��MOVB RADAPT_INERP ��FRIC�
C�OL_P M�
G�RAV��� HI9S��DSP?��HIFT_ERR-O�  �NAp�MCHY SwAR�M_PARA#� d7ANGC zM2pCLDE��CALIB� D~B$GEAR�=2� RING���<$1_8k � �FMS*�t *v M_LIF��u,(8*���M(DSTB0+_0>*_���*#z&+�CL_TIM�P�CCOMi�FB�k M� �MAL_F�EC�S�P!�Q%XO $3PS� �TI���%��"r $DTY�?R. l*1END�14�$1�ACT1T#4V22\93\94\9�5\96\6_OVR\6� GA[7�2h7�2�u7�2�7�2�7�2�8F�RMZ\6DE�D=X\6CURL� HSZ27Fh1DGu1DG��1DG�1DG�1DCNA�!1?( �PLܪ + ��ST}A23TRQ_M�d�/@K"�FSX�JUY�JZ�II�JI�J�I�E�$U1SS ? ���6Q�����+PVERS�I� 4W � �:�$' �1 TX } �� 	 ���_�_�_�U��l-�� �	������ w� ��_�_o o 9o$j_P��Ym)eAQ�o�ol����������������� �5no�ojo�l�o�o�85p����-��� :��.x �dx�fBB�!}p B |p ��p�p: ��G��<7 *�����·D�ߔ ���m�k��n�׬����.��Q ����d��o��)���=L̙�4�[�?�\���@�|�����ŏ׏������1�C�U�g�� �6U��������:T  2����'�9�@K�]�o�������<�� ��ϯ����)�;��M�_�q�����7P���$$ 1q\��aIr��Hu��H3��K����K*,*I)��mM��O��5<O$��I��{�I 3IW��ξmBo��|�B�hmz�8IB�$(�A�����ak��Lo�o�d�z� No�i�P|��P	 p�Jt�JpZ�wJ��*�/6���6S�Ir�CH�u�sH3�KK���	Ӱ2I)=j��T�{�_�ߠ[�8�#�\���{����� c{�Q� T�E��й������ݯ����F�����4T���zT���T����T��DT����T���T�{��T�vST�y�X�����T���T��gS�|P ��  ��V�	�?P�o��%����%���%����%���&��C㮈�&����&�O���K�-���"����������$���ԁ@���9�״t)w�-�����������t��ig��u��f��]�y�O� ��� �;�57�����@���? `6�� � �� Ki �����\��\���\��\��SZZ���]}�YsY�� 0�} O��G��X�Y��ѫ��r� �~n �t>� ˉt �(�� ˇo����������A����������K�E?�JT�˿���˾� xE� �
�����3����T������� k�� f�� _�*Es��+�4����4��4�2��4�g�4�����4�5�Y��5���h����_����-���6߮�� (������������$����
���~�� ��\� �`o ��a� ��� �����0 �ݞ� �� ��� �� ���� ��� ��� �I���� 
�� �,� � ��� K #��/=
dO
��O2OR(�����fe�Z�;���7�������_U����� �{�Xb���bhA���DP����k�������Ya��BR>T7P�7P0��7P�7P�/z�)*�D04�'�VՈAQ�	�	ퟱ�N龫�i�����%��h'����
�������\�����7P�  x7P��	��X��or+#00?������9���>f'xw/�- ȗ'�%�"ek}�/�/�/���m	'j!?3? '��(��+���Q�Q�G4*c4�@ @�@gs0@?�@7�@
}H�4}@%�0���9�`�8��@�r�Y@�߲@+w�0">��j�?}H�?���?���0�ī�?@��?@��c?@� ?@��M??% �3�K?>R{?>5���Ö�����>�?;���?
��?
��[�pʿUr���M�l�R�j@m�Ѿ�y�����$���`���Vž���+C�Ͼ�����L?��O����>�Nd���>��9O@�?^A?0��?7]�?4��_AB|q5�|���|�����|�����C��M��oq��a�|=Ԛl=˗�ܼ��3�|}��;��;��B���s?2�??��=�A�ѿ����������ӿ��ʿ��1�C�ֆ��:����S_�E��J�nC��ǿ��oȿ���@����̿��V���%d��Sl�Pf�BL8��L�)Pe�K�X�J��'S���M&��M5f���;��Z��U��I�6�����KQ�,����8���o�Ͽ�a[Q{�,(�$S108_PK?_T50N8Z |_ ��k_�_�_�_�_�_o �_�_oo\oCoUogo�yo�o�o�o�l2_DR_T46N6�o��m4�e�n9�bC?OMUM35=�j�6�c2�on|POU�NCE_STA7������sRpP�ROC1���`PICK
��.�k�R����v���ŏ���$P�LCL��ҕ?� nQ�?���S�6�O�Z� E�~�i�������؟ß ��� �2�