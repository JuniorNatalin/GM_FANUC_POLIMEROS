��   F�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ��	��SLGN_SET�UP_T  �H HPROC_�WET_RUN � UIF_CYCLE_TIF =JLASTMV?GUN_ON1 W	�n VVOLUME�V
� VSEAL_�AMO YATOM_AIRV�PRESSUR1��2VPART_�IDF JOB_CST�T�n^ �:�n����E�e��� � S ��SCHwEDUQ NUM��TASK�FIN�IS�F�C NI�NGFSLS.W�IZ� SLCS�TM_CTR���LOe�TPP��BFRCALL���G�DSB_�AP_# FDEFAULT_AC��JNTWARN_�EN,"USENO?NE4MAIE� {_F6 INTF��MAJb*SEQ_�IMPv*_!g%RE�COV�OK|7�60�AD�MC{SD�,REFC���"S� Ef!4�*5��*6�*7�*8�*9�*10-;�08�08�3-;�+1�+1;1P; .:,;2;8R�  ��7��7h1�8�!�8|�!�4SHORT��!H�0DUBYTE�AH�PIh1PI��!& PL_R_�EL11 @ �I��"ATA_�TYPk�BIND�EX�VAR� Rf�=�$J2$�G�21�O�O�O�H��H�C,$ R�� f!_ARY �2 ;Q�1BT� PL, SPR_R0�^X�_W�2 ^XB^XB^X1mY1 mY1mY,1mX:2�Yi\ X2�Y�\v2�Y�\�2�Y@�\�2�Y�\�2mWIhR�hY2�hh2�h�"�h �"�h2�h2�h2�h ,2�g:3.x�lX3.x�l v3.x�l�3.x	|�3.x()|�3^VBhR�x� �yh1�y�!�y�!�y1 �y1�y1�y,1�x:2 m��|X2m�	�v2m�)� �2m�I��2m�i��2�wShQ%�� ,�h0 ,�� ,�� ,�0,�0 ,�0,�,0,�:1��)� X1��I�v1��i��1������1�����1%���,T �P�OSSIBQ OP�T }!LECT�EDz�� EQUI�0 �DM_FACT�O�IDQ FLO�WCM���_BIASV� ��� ��oPURG�0AT���n ǡ0Ih1PU_P�DTH|�!�>k#X_WAI�#ISP_SIG;��_!C�ån T� Y�2�Z�S�"R�����_�Cj"HI�*�L�O��VC3�����INù4��̳�3�� �α��������� �k"�9���29�XŮC�MOD�c�L�N_
 y�TMOU�_!��GRAVI�TEP C�+�_!Sࡨ4ą����_CNpu���â�_SQ� �  ġ
��L0Y!�)֢�A2(�F� ���3���3���3��C ��C���R���R���R ���Rb��Rb�j�cb� ��8cY�j�ġw�ġ�� ġ��ġ��ġ��ġ ��ġ������#���0�9�8c
 2P@PH$���SPEED1i_����2��NOΰ�a�P��R )�EPA �R������2��B���W���A��O�G�Ŏ_��VHOȄ: �A%飚�SAMPQ ����
 ���_O -AF^�S_D0S -A3��_N{��N�LOO�����BER��CON�Vc�)+�IO_C�OU��LDBGF�L�X�cRC_D�ELA��BRA�KEu�OVRL~"TBF_OFS	T`�S^��kO �MOPGGC�URR�Zz�AU�TO_�_T{F�DU����FZ �%̡AN � ��PcRP. �.OC6�|u�q OC_LA�mO�REe�THG �A��{ �T1V�A`w������SM� FP���H _����<O �DJDL��
 4����������������%����SEC�D���PR��BI J�cZ&2�Z&�2Z&B�Z%2c*2q*2*2R�x�2��%`�����!Hw1F�d�62�6 �26R�	5B6�R6 �R6�R6�R7�R7 ;c7-;8cF���4 55��4�9I5V��4e5 l��4�5���5�9�6�� �5;4����~CĥڣA ָ2��5?LPu�F�7���Ey��DRM�T�@�����BU�BT���� _OL�D_IS��)REQ� ��C��_ST=A��  IQW��9"TYPPRB;�CcOM��DU+ЉU ���@�XN�U�� �$� N�� �#��m�VYr�Vir�V yr�V�r�V�r�V�r�V�r�#R`�j�Efw��'�j��2��UBYTEj��h2�iiq�i�yq�(�SL�PL_P_��i� \ J��� g86���RAM�e�b 3s |Yswir�cQQi��� _�aLAz�R��2 ���_NA��%EX�JP+�FAUL��BOOKMARK��N��TCPF�LS"】w����x�v�?RTD�P�s�w����D���u�w���x���MQBIT�m*�f��w���K����AVG��TOe�������� C��_m���R���R���b��bIQJa�� ��2���B�������I2N�TR�R0T�@�2� ?�B�?���?�:�W2?� e2?�s2?��2?���Ϙ�J���Ϙj��Ϙ:�1���1��1��1ʜ2ڛII��Q��s���R �b�b�#b�1b �?b��1������� �������ʬ9��@�Y��
�y���BI����aιB�ι�aι I1ιW1ιe1ιs1ι�1θ��ηSI���`� �`m�B�mʽ`m�I0m� W0m�e0m�s0mʁ0m����% ��S|6�:u � 	�pMQON q<PLR��t����%Յ��Q_E8�$�U�wU7�o�rv�?�ATUDP { �`USRC� � � �CUSX��AFLO�W_CMN�FL^��D_TY����ID���н�ACC�����S �����IN�@�Кs��%���@2��Q-��7�ND� �}�5��P�D�Й���հ����_�_�_�BoTo�B���" ���$$CpS � ���L� �  T� A�V�ERSIONI��  �:o�$SL� EQI�lT�u� r����{�EQ
!��X�q���{�GNS�Q2 j���,����T�*����	-�9SLWIZARD9f��� ������{�S�2���  �sT�CT�)?���(@�{d  ����2�^A ~jE� C�^� �� =������� �///�(H%�H) H/f'/�/�/>/l/b/ t/�/?!?�/�/<?"?X{?�?s�T��,��?n(MOV_HOlp�?�8�3Q�?��?Р�7OEJ@ 5@T���CH!m@g  S�EH{���T�
EM��?�O�O�I�EB�3~�?�1�T��34PNT �O;_2�<P]0?B?�_�b_�_�_�?n�_q3 �/,k�T��~��  '�P,i=,oro�o�oYo �o�o�o�o&8 �o\n�C��� �So�
��.��R� d�v�9�������Џ�� ���ۏ<�N�`�r� ��������̟ޟ�� �&�8�J�V�%V�z� e�����¯���ѯ
� ��@�+�d�O���s� �������Ϳ��*� �N�9�rτ�oϨϓ� �Ϸ��������&�J� 5�n��L�ߡ߳�X� 0B���_x5�Y� ������/����/ |_r_�/1�C�U���� p�&�����h_����^? -?�?�?��?�  O�$O�HOZOlO~O �O�_q}��O�_  _�D_���4/�_ [/m/���/
oo.o @o�?!?3?E??i? {?�?P?�?�?�?�?�? OO/O�?SOeOwO� HO�O�O�O�O�O__ +_�OO_a_s_6_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�o�o�o�o �o�o�o^�#G2 kV������ ���1��U�g�R� ��v�����ӏ����	� �-��Q�<�u�`��� ����ϟ���ޟ���;�M�_�  �$S�LSTATUS �2������� b��� ��ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�w� � #�Ϸ���������� #�5�G�Y�k�}ߏߡ� ������������
� C�.�g�R��v��� ������	���-��Q� <�u������������� ��);M_q ������� %7I[mf� ������/!/ 3/E/W/i/{/�/�/�/ �/�/�/�/�??A? ,?e?w?b?�?�?�?�? �?�?O�?+O=O(OaO�LO�Oj�USRCSoT 2�� X�F	�H�E�O�J�O_� _2_D_V_m�VOLSET1  0�OG�O�mZ2{_�nY3�_nY4�_nY5�_  