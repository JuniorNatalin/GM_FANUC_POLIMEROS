��   @�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����SEAL_MAP�_T  0 ��DI_��_RD�YT 8ICF�LTB	] QDIS�P>	wQFULL�OPNB��	CL�S�	� �LT_S�TRB��QPRSSRRMB�Q`� �BQHI8/Q( SELBN�QVOL�
ko	ESTP	�o
]��QCOM��QB�UBL\	�oRM�1EMT~$(2�,."QMATW�BK$C)HIR)HI~C&TR_EMP_�%}(N�,�"})��)�o
MOD
� o	�NSNG		1	W0j'2'GH(9C5~QNOT_CASc4�&0RA_�5�?ART_OK��36QIN� OCB�4C'J\	�4C&�0�9�3�c�7CQAUTO�)5EC'NU�)UEo?EPRESE�'vD�'UM+�CQ� I�N�0B�E�DETE�6�E})� \G�D�ICHKP�U[�Fn&5U�R_AD�V�VT�URGRQUE�vTmY�A}Y��A�HG_BRSqH��Ty8_BYW�UQ�0E1B�R�ZU2�Z2�Z3�Z3�ZU4�Z4�Z5�Z5QG�NU�~gye�P_AC�3�gyew)5 �hye�X�fQAiw B�g�eK!�  ut{ c2w�e�XPvKz;vi?O_ONGU��t �zd�u�z2d�u�zNd��u�zjd�u�z6�z6 �wuQ|T/�)��xQ�)� �xq�)��x��)��x�� )��у�u�P�톃u�] ���uAB��EqQ�u+��uSET(7�G��ukC� `��uCL� ^��A�� � P����uRLD�����G_W�0؛�ut�T �����v�A�) Q;�~�uEND_JO��]��uGOO_�{�熇ANE@�v����F
��F��M���ۥ�u w��u���vB��p��;��uWAIqn$W�#�DVTR2�z��vKTOuQ�v��}�8�����uBLK��ٵ��uUTH����ѶS ���󩈙�7�h0A�<h0)�INCH�y� q�V���A��X�űʪv }{-i�ű��vWi���v�si�_I�#B�=�RAl�^�=��i��v�c���c��MD�1 s��~��ATM_AI��ש�w@�t����S�SUR|S
��HA�N��;t+��Sy��$��$$CLASS  ���r�j��!��!g�VE+p�ONo� � �:�$SL�IO,  2 ��!� ������ ���������	��D� V���z���w������������
��q�+Rs�(��� ��� DV 9z�����_H�
/-	/,
B, 9/+u/�/q/�/�/�/ �/�/?�/�/B?-?f? x?�?�?�?�?�?M?�? QO,O>O�[OmO� �O�O�O�O�O�O_�O (_:_L_^_p_�_�_O !_�_%/�_I/�_�6