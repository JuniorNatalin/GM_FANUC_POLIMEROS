��   ��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����PMC_CFG_�T   � �$'NUM_MS�K  $EX�E_TYPECM�EM_OPTPN�_CNFCIF_�CY:gSCN_�TIME E R?ESET_P�D�o LJ �HECK�_DSBLC $�DRA> ARGI=NCSTORJ���&DEV. d� 	7OC'HA�R�ADD�SI�ZORACBSLmO[ODKIOKOCCPYC&l >/  L ��ph99IDX��&L. � �
�EQPLHR�AT�TRKBU�F| ��UN_�STATUS�C�U��MAX(I���SNP_PA��  � �� ANNE�� O~W CTION_��PU�   �$BAUD�N�OISYmN�T�1�#2�#3�$_P�R�T4P' DA�TA�CQUEU�E� PTH[$MM�_��%&!RETR�IESCAUTOb!R[��BG �� �ISP_IN�Fd�' CLIM9I� B5AD_H C3 H��#d6�#d6�#d6 �#W1� �#�4�#�4�#��4�" ��$$�CLASS  O����1����=�0VERSg �8��0�:��iFG0 �5���
@+A�2������d��3CC�  2uG'@d $)D xO��uO�O�O�O�O�O �O__:_)_^_M_�_ q_�_�_�_�_�_�_o o6o%oZoIo~omo�o �o�o�o�o�o�o2 !VEzi��� ���
��.��R� A�v�e���������� я���*��N�=�r� a���������ޟ͟� �&��J�9�n�]��� ������گɯ���"� �F�5�j�Y���}��� ��ֿſ�����B� 1�f�Uϊ�yϮϝ��� �������	�>�-�b� Q߆�uߪߙ��߽��� ����:�)�^�M�� q����������� �6�%�Z�I�~�m��� ������������2 !VEzi��� ���
�.R Ave����� �/�*//N/=/R,�CIF 2aKP+ )DX5D�)G�&UȪ'�%Y�(�(��!�%� �&D6C�>9@  '^/X/ "?K?F?X?j?�?�?�? �?�?�?�?�?#OO0O BOkOfOxO�O�O�O�O �O�O�O__C_>_P_ b_�_�_�_�_�_�_�_ �_oo(o:oco^opo �o�o�o�o�o�o�o  ;6HZ�~� ������� � 2�[�V�h�z������� ����
�3�.�@� R�{�v�����ß��П����#TYPE �2�+ (�#5	0d�����!����h���	0��ɯ	0������~#SNP_PA?RAM �+���1'C�q�ꦠ�!ۤ�"��1	0U D��)R�