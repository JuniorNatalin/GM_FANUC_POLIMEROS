��   F�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ��	��SLGN_SET�UP_T  �H HPROC_�WET_RUN � UIF_CYCLE_TIF =JLASTMV?GUN_ON1 W	�n VVOLUME�V
� VSEAL_�AMO YATOM_AIRV�PRESSUR1��2VPART_�IDF JOB_CST�T�n^ �:�n����E�e��� � S ��SCHwEDUQ NUM��TASK�FIN�IS�F�C NI�NGFSLS.W�IZ� SLCS�TM_CTR���LOe�TPP��BFRCALL���G�DSB_�AP_# FDEFAULT_AC��JNTWARN_�EN,"USENO?NE4MAIE� {_F6 INTF��MAJb*SEQ_�IMPv*_!g%RE�COV�OK|7�60�AD�MC{SD�,REFC���"S� Ef!4�*5��*6�*7�*8�*9�*10-;�08�08�3-;�+1�+1;1P; .:,;2;8R�  ��7��7h1�8�!�8|�!�4SHORT��!H�0DUBYTE�AH�PIh1PI��!& PL_R_�EL11 @ �I��"ATA_�TYPk�BIND�EX�VAR� Rf�=�$J2 d�G21�O�O�O�O+�$ R� f!_�ARY 2 �;Q�1BT P�L, SPR_R0 �^X�_W�2^XB^X B^X1mY1mY1mY ,1mX:2�Yi\X2�Y�\ v2�Y�\�2�Y�\�2�Y(�\�2mWIhR�hY2 �hh2�h�"�h�"�h2 �h2�h2�h,2�g:3 .x�lX3.x�lv3.x�l �3.x	|�3.x)|�3^VBhR�x��yh1�y �!�y�!�y1�y1�y 1�y,1�x:2m��|X2 m�	�v2m�)��2m�I���2m�i��2�wShQ%�� ,�h0,�� ,� � ,�0,�0,�0,� ,0,�:1��)�X1��I� v1��i��1�����1������1%��,�T �POSS�IBQ OPT ~}!LECTEDz��� EQUI0 �DM�_FACTO�I�DQ FLOWCM����_BIAS�V� ��� ��PURG�0AT��n ǡ�0Ih1PU_P�D�TH|�!�k#X_�WAI�#ISP_SIG;�_!C�åRn T� Y�2Z�S�"�R�����_Cj"H�I�*�LO��V1C3�����INù4� �̳�3���α�� ��������k"��9���29�X�C�MOuD�c�LN_
 y�TMOU_!�ĿGRAVITEP C�+�_!S��4ą����_CNu����_SQ�   ġ
��LY!�)���A2(�F����3�� �3���3��C��C�� �R���R���R���Rb� �Rb�j�cbք�8cY� j�ġw�ġ��ġ�� ġ��ġ��ġ��ġ�� ����#����9�8c�
 2P@PH$��S?PEED1_����M2��NOΰa�P��R )�EPA�R�� ����2�B���4W���A��OG�Ŏ_��VHO�: Qy%飚�SAMPQ  ����
 ��_O -AF^�S_DS -A3�Ɛ_N{���LO�O����BER>��CONVc�)~+�IO_COU��?LDBGFL�X��cRC_DELA~��BRAKEuހOVRL"TB/F_OFST`�aS^��kO MOP�GGCURR��Zz�AUTO_��_T{�DUh����FZ %̡qAN � ��PRP.� �.OC6�u�q O�C_LA�O�R-Ee�THG A��{ �T1V�Aw���,���SM� FP��тH _����O �D'JDL��
 4���� �����������%<����SECD���PR��BIJ�cZ&@2�Z&�2Z&BZ%2c*�2q*2*2R�x�2���%`�����!Hw1 F�d�62�6�26R� 	5B6�R6�R6�R 6�R7�R7;c7 -;8cF���455��4 �9I5V��4e5l��4�5 ���5�9�6���5;4�� ��~CĥڣAָ2��5?LPuF�7��8�Ey��DRMT�@��x���BUBT����� _OLD_IS��)REQ ���C��_STA�� � IQW�9"TYvPPRB;�COM����DU�+ЉU Д��@�XN�U� �$� N���#��m �VYr�Vir�Vyr�V�r��V�r�V�r�V�r�#R `�j�Efw��'j��2��UBYTEj���h2�iiq�iyq �"��SLPL_�P_��i� \ J��� g6���RAM�e�b3s |Ys�wir�cQQi��[ _�aLA�R���2 ��_NA���%EXJP+�F�AUL��BOOK�MARK����TC	PF�LS"�w����x�v�?RT�P�s�w����D���u�w��p�x���MQBIT� m*�f��w��K�����AVG��TO�e�������� C��_ m���R���R��b��bIQJa����2���@B�������I2N�TR�R0T�@�2�?�B�?� ��?�:�W2?�e2?�s2 ?��2?���ϘJ���ϘPj��Ϙ:�1��1��U1��1ʜ2ڛII� �Q��s���R�b� b�#b�1b�?b� �1������������ ��ʬ9���Y��(
�y���BI����a ιB�ι�aιI1ιW1 ιe1ιs1ι�1θ��ηSI���`ǝ`m�B� mʽ`m�I0m�W0m�e0�m�s0mʁ0m���%� 4�S6�:u� � 	�pMQON  q<PLR�t����8%Յ��Q_E8�$��U�wU7�o�rv?�AT�UDP 7�aU�SRC� w� � CUSX���AFLOW_CM�N�FL��D_T5Y���ID����.��ACC�����0S �����IN�@�� �s��%���2��Q-��7�ND�}�5��P�D�Й���հ� ���_�_�_BoTo�B����" ��$$�CpS  �{��L�   T�� A�VERSI�ONI� � �:�$SL�� EQI�T�u� fr����{�EQ
!Ѕ�X�q��{�GN�S�Q2 j���q,����T�*�����	-9SLWIZARD9 f����������{�S2����  �sT�C�T�)?��(@��{d  ���2��^A jE�g C�^� ��� =��� �����///� (H%�H)H/f'/�/ �/>/l/b/t/�/?!?��/�/<?"?{?�?s��T��,�?n(?MOV_HOlp�? �8�3Q�?�?Р�7OZEJ@ @T���sCH!m@  S�VEH{���T�
EM���?�O�O�I�EBP�3~�?�1T��34PNT�O;_2�< P]0?B?�_b_�_�_�?8n�_q �/,k��T���� W '�P,i=,o ro�o�oYo�o�o�o�o &8�o\n� C����So�
� �.��R�d�v�9��� ����Џ�����ۏ <�N�`�r��������� ̟ޟ���&�8�J�V�%V�z�e�����¯ ���ѯ
���@�+� d�O���s�������� Ϳ��*��N�9�r� ��oϨϓ��Ϸ����� ���&�J�5�n��L���߱���0B�� �_x5�Y����� ���/����/|_r_�/ 1�C�U����p�&��� ��h_����^?-? �?�?��?� O�$O �HOZOlO~O�O�_ q}��O�_ _�D_ ���4/�_[/m/�� �/
oo.o@o�? !?3?E??i?{?�?P? �?�?�?�?�?OO/O �?SOeOwO�HO�O�O �O�O�O__+_�OO_ a_s_6_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o ^�#G2kV� �������� 1��U�g�R���v��� ��ӏ����	��-�� Q�<�u�`�������ϟ ���ޟ��;�M�_��  �$SLST�ATUS 2�������� �ԗ��� ��ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/� A�S�e�w� �#�Ϸ� ���������#�5�G� Y�k�}ߏߡ߳����� ������
�C�.�g� R��v��������� 	���-��Q�<�u��� ������������ );M_q��� ����%7 I[mf���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/�??A?,?e?w? b?�?�?�?�?�?�?O �?+O=O(OaOLO�Oj��USRCST 2-�� X�F�H�E�O�J�O_ _2_D_�V_m�VOLSET�1  0�G�OI�mZ2{_nY3�_�nY4�_nY5�_  