��   �i�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DCSS_CPC�_T   � �$COMMEN�T $EN�ABLE 6 M�ODJGRP_N�UMKL\  $UFRM\~] _VTX 6 ~�   $Y�{Z1K $Z2��STOP_TYP�KDSBIO�I�DXKENBL_�CALMD�US�E_PREDIC�?  &S. Ǆ 8J\TC��u
SPD_LI`_���SOL��&Y0  � �1CHG_SIZ�$APGE.SDIS��GB�C����J
p 	�J�� &��"�))$'2_SyE�� XPANI�N��STA�T/ D $�FP_BASE �$_ K�$!Y �&_V�.H�#� �&J- q�ZAXS\7UPRJLW7S<e� ��$� | 
�/�/�/�D&?8?z�&EL�EM/ T ��2�"NOG�0�3�UTOOi�2HA�D�� $DAT=A" �&e�0  @@p:�0 _2 
&Pp%' � p!U*n   �FS�Cz�B�� �B(�F�D(�R|UC�DROBOT�H��CqBo�E�F$OCUR_2R &�SETU�	 l|� �P_MGN�INP_ASS� 0"@�� �3�8B7gP@@U�^V�Sp!��&T1�
`B|8�8�TM 0 6P�+ Ke�1VRFY�8
dD5F1�� ��W��1k$R��&TPH/ ({ �CA�CAt�CA3�BOX/ 8�0����У�b'oEc��TUI}R�0  ,{ �FR`ER�02 {$�` �a�_S�b(�fZN>/ 0 {9F02� -a0rZ_0��_0�u0  @�Q�Yv	�o:n���$$CLLP  O����q��Q���Q�pVERSIO�N�x  ��:�$' 2� �xQ   ��!A CART? 50_60���p� �p�q����8��Z� ��A���1�Ö � �;�M�����/� Da��
�� ���pool cart 70_8
�|�.�m� �Th�~V�E@ �H� z���2 ���qF���ŉ S�;�W�􏕟��͟<� �`�r�����(�]�o� ޟ����J�ۯʯ������Fence By C������>яg@ �z����/�����*�by Gate=�O�a�O]� ė���E?��A� �E@Hϛ�
�ݱ 0�c��� �w�E@�.�g����ϖ�0�Stairs Low����3�C�<���l�;�ADw����Ϙ�ݏhigh0�B�4�D��E�u߇����C����Զ%�corner������_�C��+����B_���fյplatform�χ�1���w��U�ŧ���u� ����conve�yoy��)�;�b�E5t�����r���ߙ��0�etween�������>��T�^�C���/�b�D�υ�� �����5j|� �!W��// �B/����/��/ �///�/S/e/w/,?�/ P?b?�/�?�/??�? =?�?Os?(O:O�?�? pO�?�O�OO'O�OKO ]O_�O6_H_Z_�O~_ �O�O�_#_�_�_�_k_  o�_�_Vo�_zo�o�o o�o1oCoyogo�o. @�od�o�o�� ��Q�u��N� �r�������)�;� ��_��&���J���ˏ ݏ�����ȟ7���� m��4���X�j�ٟ� ���!�֯E����� ��B���ïx�篜��� ��/��S�e�ω�>��P�b�i�$DCS�S_CSC 2�{ ��Q  Dֿ��~*� ���ϼ���#���5�� k�:ߏ�^߳߂��ߦ� �������C��$�y� H��l�������	� ��-���Q� �2���V� ��z����������� ;
_.@��v�	�z�GRP 2N�� ���	<� !E0iT�x �����/�// /S/>/w/b/�/�/�/ �/�/�/�/??=?(? a?L?�?�?�?t?�?�? �?O�?'OOKO6OoO �O�O^O�O�O�O�O�O _�O5_ _Y_k_}_H_ �_�_�_�_�_�_�_o 
oCoUogo2o�ovo�o �o�o�o�o	�o-? Qu`����������_GS?TAT 2����,8��b��>�5�R��>���?b�f�:�y2==�=Ǽ�������	��D�?a&D�fۇ���8V�d��>�����v8����)?�  ��?���4��ZË\�C2����V����ga>nӤ�?Z�4?C{)��ħ0?�K����BK�C�u��De�ƅ>v������?v��ʾ�Ö������(?\E1��ݗ.���?��4�oC����D��8��u�x���Pv���/�"�7&�>�;?�d�n9ׯ���
:�D��D���ƅ�da�>�Ӂ�R����W��[��ׅ���==�<��t?{�c�Y�k�}����� ������(�:��^� p�����	ɒ��ƅ�� ̯��ȯ���� �"� 4�V���j�����ćv� �B��&�8��\�n� ��¿�Ϟ����ϸ��� ����:�$�F�p�Z� lߦߐ�N���������0��T�f�D�b��>�'�T���>�����*:����=>�����/�����	�D�f9D�P����J>��䞃w�����֪�䲀J���C�4o�>n�ޔ?Z�??C�x�ĦR?��+���BO�C�|$De�6������,�?v����ۖ�L�����?\K9��ݟƾ�����4мC��A�D��x6�~-�W���:�J�7N���R�>�!S?d���9���
�?tD�,D���n�_O>�Կ]�T���������ڛ�>�?�<�.|?��� ����J�.R dB���Ϻ���� ���0,f Pb�����z /&/xJ/\/:/�/�/ ���/��/�/�/�/ ??$?F?p?Z?|?�? �?�?�?/OOp/BO TO2OdO�OhO������ ����������(�:� L�^�p����������� �O�O �OLo�O<o�o �oro�o�o�/�?�o�?  *6`Jl� ��������o D�V�4�z���j��� �o�����"��.� X�B�T���x������� ������<�N���r� ��b������O
oo�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ ���0oj�|ϖ��ϲ� ������Ώ���$��� 0�Z�D�fߐ�zߜ��� ���������2���� t���d�������� �F��"�(�R�<�^� ��r������������� ��*��l~\� ����ԯ:�L�
� �.�@�R�d�v����� ����п����� &`Ϛ/�/��/�/ �/??��(B?L>? `?b?t?�?�?�?�?�? �?O,OO8ObOT�O �O�/�O�O�O�O_*? <?vOL_ROX_�_l_�_ �_�_�_�_�_�_$oo 0oZoDo"_�o�O�o�o �o�oX/j/|/: L^p����� �� /J/$/6/H/2 DV�oʏ܏�� �� ��6�H�._hor�|o~� ������ޟȟڟ���� �2�\�F�h����o¯ ԯ&���
��.�@�Z� ��j���f��������� �ҿ����*�T�>� `ϊϰ��������� ���8�߈�����j |������� ��0�B�T�f�l�b� t߮�(������0�B�  �f�x�^��Ϣ�tϮ� ��������D. @zdv��X�� �(:^p�� �������/ �/$/&/8/Z/�/n/ �/�/��/�/N ?2? ?V?h?R߸���ߚ� �߾���������*� <�N�`�r����? �?��x?*_|?:_`_>_ P_�_�_��/�_�/�_ o�_o>o(oJoto^o �o�o�o�o�o�o�_" 4XjH���_ �o��o� ���6�  �B�l�V�h������� ����,�
�P�b��@������u�$DC�SS_JPC 2��uQ ( D���������0ԟ)���
� _�.�@�R���v����� ﯾ���7���Z� �N�`����������� ̿!��E��i�8ύ� \�n��ϒϤ϶���� ���S�"�w�Fߛ�j� |߾��߲�������� �a�0��T��x��� ��������'����� o�>�}�b��������� ������"G(} L^p���� �1 U$6�Z l~����/� ?//c/2/D/�/�/z/ �/�/�/�/�/)?�/M? ?q?@?�?d?�?�?�? �?�?�?�?7OOEO�*��S��Ý@0O�O TO&O�O�O�O�O!_�O _W_*_<_N_�_r_�_ �_�_�_�_o�_o@o eo8oJo�ono�o�o�o �o�o�o'a4 F�j|���� ����]�0�B��� ��x���ۏ����ҏ#� ���Y�,�g�P���t� ��ן����Ο��� U�(�:�L���p����� 寸�ʯ��?��c� 6�H���l�����ῴ� ƿ�����_�2�D� ��h�zό��ϰ��� � %���
�[�.��Rߣ� v߈��߬�����!�����W�*�<�pHMOD�EL 2�K�xTool �CHANGE��
� <v�cz����C�K���  ��m� C�  "��D��K�����I� ����E��'�t�K�]� ��������������( ��^5GY�} ����M���� �p�Yk}� ����$/�// 1/C/U/�/y/�/�/�/ �/�/�/�/	?V?-??? �?'9g?y?�?a?�? �?.OOOdO;OMO�O qO�O�O�O�O�O_�O _N_%_7_I_�_m__ �_�_�_o�?�?�?�_ o�_EoWo�o{o�o�o �o�o�o�o�oX/ A�ew���� ���B��+�=�o ��7oe�w�M���͏� ��P�'�9�K�]�o� ��Ο�����۟��� �#�5���Y�k����� ���������ۯ�Z� 1�C���g�y�ƿ���� ������D��-�z� Q�c�u��ϙϫ����� ��.���)�����#� Q�c��ߧ߹������ ��%�7��[�m�� ����������8�� !�n�E�W�i�{����� u���������F/ |Sew���� ��0+=O a������� �//��t/=/O/ �/�/�/�/�/�/�/:? ?#?p?G?Y?�?}?�? �?�?�?�?$O�?OZO 1OCOUO�OyO�Oa/s/ �/�O�O2_�O_-_?_ Q_c_�_�_�_�_�_�_ �_�_oodo;oMo�o qo�o�o�o�o�o�o N�O�O);�# �����&��� \�3�E�W�i�{���ڏ ��Ï������/� A���e�w�ğ_q�� �������f�=�O� ��s���ү����ͯ� ��P�'�9���]�o� ��ο�����ۿ�:� ՟���'�9��}Ϗ� �ϳ���������� 1�Cߐ�g�y��ߝ߯� ��������D��-�z� Q�c�u�K���oϝ�� �����R�)�;���_� q������������� <%7I[m� ��������J ��%�i{�� �����F//// |/S/e/�/�/�/�/�/ �/�/0???f?=?O? a?7�?[�?�?O�? �?>OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_p_G_Y_�_}_�_�_�_�_�_�:�$D�CSS_PSTA�T ����AaQ    �6�T``l  bn(`to�o�o�odo �k  `B`�ar`o$�9cAeN�`C�u~2dSETUP ;	AiB�dZd��1�t-iT1SC �2
�z�`�1Cz�3����uCP [R�|��0D�? X�j��?��������֏ ���ɏ�0�B��f� x�G������������ �ן,�>�P��t��� ��g���ί�>F��� ��9�K�]�,������� t�ɿۿ���#�� �Y�k�:Ϗϡϳς� ���������1�C�� g�y������H��� ��	���-�?�Q� �u� ���h������� ���;�M�_�.����� ��v���������% �ߞ�[m����� �����!3E i{J\��� ��/�//A/S/"/ w/�/�/j/�/�/8J ??�/=?O?a?0?�? �?�?x?�?�?�?�?O 'O�?O]OoO>O�O�O �O�O�O�O�O�O#_5_ G__k_}_�/�/�_�_ L_�_�_o�_1oCoUo $oyo�o�olo�o�o�o �o	�o?Qc2 ���z���� �)��_�__�q���� ������ݏ��Џ%� 7�I��m��N�`��� ǟ������ޟ3�E� W�&�{�����n�ïկ <�N�����A�S�e� 4�������|�ѿ��� Ŀ�+����a�s�B� �ϩϻϊ�������π'�9�K��o߁ߑ���$DCSS_TC�PMAP  ������Q_ @ \�\Х\�\���\��\�\�\�	�� � \�\�\��\�\�\�\��\�\�\�\�J\�\�\�\�\�U\�\�\�\�U\� \�!\�"\�U#\�$\�%\�&\�U'\�(\�)\�*\�U+\�,\�-\�.\�U/\�0\�1\�2\�U3\�4\�5\�6\�U7\�8\�9\�:\�U;\�<\�=\�>\��?\�@��UIROw 2�������� ��$�6�H� Z�l�~�����������@���� 2[��� [������� ��!3EWi {���<�`� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?�a?��?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O�T?�O��UIZN �2��	 ��� ��._@_R_W�)_~_�_ �_e_�_�_�_�_o o 2o�_VohozoIo�o�o �o�o�o�o
�o.@ Rd'��i{� ����*�<��`� r���G�����̏���� ��׏8�J�\�+��� ������y�ڟ쟻���"�4��O��UFRM� R�����8 _ߌ���]�¯ԯ���� 
��.�@��d�v�Q� ������п⿽��� �)�N�`�w��ϖ�5� ���ϧ������&�8� �\�n�Iߒߤ�ߵ� �������"���F�X� o�|��-������� �����0��A�f�x� S������������� ��>Pg�t�% ������( :^pK��� ��� //�6/H/ _V/~/�/k/�/�/�/ �/�/�/ ?2??V?h? C?�?�?y?�?�?�?�? 
O�?.O@OW/i/vO�O 'O�O�O�O�O�O�O_ *__N_`_;_�_�_q_ �_�_�_�_oo�_8o JoaOno�oo�o�o�o �o�o�o"�oFX 3i��{��� ���0�B�Yof�x� �������ҏ䏿��� �,��P�b�=����� s���Ο����ߟ(� :��