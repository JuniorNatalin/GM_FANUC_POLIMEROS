��   O�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����DMR_GRP_�T  � �$MA��R_DO�NE  $O�T_MINUS �  	GPL�N8COUNP �T REF>wPO�OtlTpBC�KLSH_SIG�oSEACHMS9T>pSPC�
��MOVB RADAPT_INERP ��FRIC�
C�OL_P M�
G�RAV��� HI9S��DSP?��HIFT_ERR-O�  �NAp�MCHY SwAR�M_PARA#� d7ANGC zM2pCLDE��CALIB� D~B$GEAR�=2� RING���<$1_8k )߀�FMS*�t *v M_LIF��u,(8*���M(DSTB0+_0>*_���*#z&+�CL_TIM�P�CCOMi�FB�k M� �MAL_F�EC�S�P!�Q%XO $3PS� �TI���%��"r $DTY�?R. l*1END�14�$1�ACT1T#4V22\93\94\9�5\96\6_OVR\6� GA[7�2h7�2�u7�2�7�2�7�2�8F�RMZ\6DE�D=X\6CURL� HSZ27Fh1DGu1DG��1DG�1DG�1DCNA�!1?( �PLܪ + ��ST}A23TRQ_M�d�/@K"�FSX�JUY�JZ�II�JI�J�I�D��$U1SS  ���6Q�����+PVER�SI� 4W  �:�$'� 1 TX � �� 	 ����_�_�_�VE0��`�������E� M��;�����_o�W��\�Q a���S�+�\c_P��TWgo?S�o�^F?� <>��6�H��P���UI�9ۈno�ojo�l�o�o�85qW������ a .w  �$�$fq��gB B �}p|p �q�p �: ��T��h"q��]��������ZV��~���A�  ~\�����T���X���d�o��)���=gL��4�[�?�\���@�|�����ŏ׏ �����1�C�U�g�� 6U��������:T  2���� '�9�K�]�o�������<����ϯ�����)�;�M�_�q�������$$ 1q\��aH?[�G���GE{�I����J�'K%���mN|��O����O}.#J���tI�B�HX�C�mBo��|���	\X)*A�Z����N���FC6%�o�d�z� O�<��P��PB���K�%J�W�I_�&�����Ϣ�S�H?^z�G��{GE��I��]Ӱ'װ�^��Ta�e_����b�Tϕieo\�a���� @P  ��B��֌ӄр� }�U��O��Q��T���S[v�S]�S]��������-��0S^,A�T,x������.���2��4��5��8���MT��T�+��SԮ ����� ���y������.�3���/����^����'����$��^º�C���G�Z�������)��*��+��,��-q3��֫�AI'>��=L;��0Ctb@����������=���@��S��S���@��@-��BqLB�Q�>��>�/����r�u�q����q6b�rQ�m�s�N�r����b�K�b��G�b��_����_l �r�����|���_���r���ro�Y�s-�sg�M�q���q��$��'W����3���b������H�B��B��'�B���Ou߿�P�C�>�H�HB����^�>���)���s��������H�������������e�������C���a7��[����S�������!ϗ�&��C�
ڜ��\����0��;����T���������������W����y����6*��\��Ը���#����<������p��V�����S~��Sp���ӣ��ӎ���"L������Z���;����Vёq�q2;
�
�;VV*	*(BR�Vd>7P��7P��S����7ߩӇ����R��e  �j����]�o ���
� 7P����.������7P�ϋ��܆��P�U'�_�7P�S�#7P�7P�7Px
7P���CR�����%7P�7P��{���s7P�BVdVl��>T
���#�� �p �7P����p5چ�=QT�7P�7PQ�(�w/�/�'�p�"�/�"���uj��/�/����"5#����o/4:=p��/O4"9"7�����#����s0�n����1�Ȥ��m~�+�� ��"���1?I���?I���0�w0(�w0Zw0�w0�s0�!��u�����п��z����迍����������1��o�7��WS��S�)���0���ž���.��������������������� !�>d�h>kt��>o:>t7��>W�s>fH��>�+�>��B�>�y�>�?�>��/A?7.�/?7�>fK�w>gU�>a���>`�E>j��8>j���2����J��	���򻯿�4����=<�ݭ�пݕ�ݷ�d��3ÿ���ăA@��?@�����;�����L�������������}�!������;�F���ҍs���2���nF��)��ŕ��Ŭ���K���H��A���7k��H9��@���Hg���O��ϧ\�ο2��@!@�)Δ@(ک@�(0h@'ɇ@�+��@)�S@���@W�@�g�@��@���+Q�K�A��K�N@)Bp�@)!�@*��@*MB@)��@(�v,($FLT_MH
?�_k_�_�_�_�_S103�_PK_TCOM�UM35_R01��_�STL_LAT�C�_
o$CUSTOOK5o6oo�olo �o�o�o�o�o�o�o�9Do]�\8PICKoj|��_�� ���7��0�m�T����x���Ǐ��PLC�L��ҕ�� D�T�?���J�~?[���S�6�O�Z�E�~� i�������؟ß���  �2�