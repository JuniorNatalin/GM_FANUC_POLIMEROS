��   h5�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����SEAL_SCH�_T  � �COMMENT� 'AMO�U= ATOM�_AIRNEQ_�ADD_DELA�YN EQUIP�dGUNONsF�FdC_FACT�OYC_BIAS�NPRE_� S_WTIMjD�EjRAMPjR�i���xS_USE�DN DUMMY.� HORM� ��SUR�FLO�W_TYP�%M�Oe jS�_OF�SMSEBRS]MGFSEM2G	2)n^ enb	n��	��GUM_D�ROP�T�$�$CLASS  ������� ��� �VERSI�ON� � �:�$SL~, ED1 2 �  d ���=/��?�E/�� m( t'j/V*+/�/�/�/s/ �/�/�/:?�/^?�/b? ?'?�?K?�?o?�?�? �?6O�?ZO�?�?O#O �OGO�O�O}O�O�O2_ D_�O_�Ok__�_�_ U_�_y_�_�_.o@o�_ o�_goo�o�o�o�o uo�o�o�o<`�o cO)�M�q� ��8��\���� %���I�ڏm������ 4�ǏE�����!��� ğW���{�럟�0�B� ՟	���i������S� ��w�篛�,�>��� ��e�Q�+������s� �Ͽ��:�Ϳ^��b� �'ϸ�K���oρϓ� ��6���Z������#� ��G��ߍ�}ߏߡ�2� D������k����� U��y����.�@��� ���g���������� u�������<`���cO) Used� in MOV_SEAM���s ��):�^�b '�K�o�� �6/�Z/��/#/ �/G/�/�/}/�/�/2? D?�/?�/k??�?�? U?�?y?�?�?.O@O�? O�?gOO�O�O�O�O uO�O�O�O<__`_�O c_O_)_�_M_�_q_�_ �_�_8o�_\o�_oo %o�oIo�omoo�o�o 4�oE�o!� �W�{��0�B� �	��i������S� ��w�珛�,�>��� ��e�Q�+�������s� �ϟ��:�͟^��b� �'���K�ܯo����� ��6�ɯZ�����#� ��G�ſ��}�����2� D�׿���k�ϰ��� Uω�y��ϝ�.�@��� ���g�߬߾ߙ߅� u����߫�<��`��� c�O�)��M���q��� ���8���\����� %���I���m������ 4��E��!� �W�{��0B �	�i��S �w��,/>/// �e/Q/+/�/�/�/s/ �/�/�/:?�/^?�/b? ?'?�?K?�?o?�?�? �?6O�?ZO�?�?O#O �OGO�O�O}O�O�O2_ D_�O_�Ok__�_�_ U_�_y_�_�_.o@o�_ o�_goo�o�o�o�o uo�o�o�o<`�o cO)�M�q� ��8��\���� %���I�ڏm������ 4�ǏE�����!��� ğW���{�럟�0�B� ՟	���i������S� ��w�篛�,�>��� ��e�Q�+������s� �Ͽ��:�Ϳ^��b� �'ϸ�K���oρϓ� ��6���Z������#� ��G��ߍ�}ߏߡ�2� D������k����� U��y����.�@��� ���g���������� u�������<`�� cO)�M�q� ��8�\� %�I�m�� 4/�E//�/!/�/ �/W/�/{/�/�/0?B? �/	?�/i??�?�?S?��?w?�?�=�$SL�SCHED2 2� ���8A  d ��? ZOO~O�?�OmO�?�O kO�O�O _�O�OV_�O z___1_C_�_g_�_ �_�_�_�_Ro�_co+o o-o?o�o�ouo�o�o 	�oN`�o'� ;��q���� J�\�7�#����o�I� ڏ��������ǏX� �|����3�E�֟i� ��������ßT��x� ��/�A�үe�㯫� ������P�b���)�� ��=�ο�s������ ��L�^��%�υ�9� ���Ϸϣϓ������ Z�5�~�߁�m�G��� k��ߏ� ����V��� z���1�C���g��� ������R���c�+� �-�?�����u����� 	��N`��'� ;��q��� J\7#�oI ����/��X/��|//�/3/E"U�sed in MOV_SEAM�/ �/�/�/?�/G/X?�/ |??�?3?E?�?i?�? �?�?�?�?TO�?xOO O/OAO�OeO�O�O�O �O�OP_b_�O)__�_ =_�_�_s_�_�_o�_ Lo^o�_%oo�o9o�o �o�o�o�o�o�oZ 5~�mG�k �� ���V��z� ��1�C�ԏg����� ������R��c�+�� -�?�П�u�����	� ��N�`��'����;� ̯ޯq��������J� \�7�#����o�I�ڿ ��������ǿX�� |�π�3�E���i��� �ϟϱ���T���x�� �/�A���e��߫ߛ� �߿�P�b���)��� =�����s������ L�^���%����9��� ������������Z 5~�mG�k �� ��V�z 1C�g�� ���R/�c/+// -/?/�/�/u/�/�/	? �/N?`?�/'??�?;? �?�?q?�?�?O�?JO \O7O#OO�OoOIO�O �O�O�O_�O�OX_�O |__�_3_E_�_i_�_ �_�_�_�_To�_xoo o/oAo�oeo�o�o�o �o�oPb�o)� =��s���� L�^��%����9�ʏ ܏��������ɏZ� 5�~����m�G�؟k� ���� ���şV��z� ��1�C�ԯg����� ������R��c�+�� -�?�п�u�����	� ��N�`��'�χ�;� ����qϥϕ�߹�J� \�7�#�߃�o�I��� ���ߑ������X��� |���3�E���i��� ������T���x�� �/�A���e������� ����Pb��)� =��s��� L^�%�9� ����/��Z/ 5/~//�/m/G/�/k/ �/�/ ?�/�/V?�/z? ??1?C?�?g?�?�? �?�?�?RO�?cO+OO -O?O�O�OuO�O�O	_ �ON_`_�O'__�_;_��_�_q_�_�_o�]��$SLSCHED�3 2 ����Va `� �_xo5o�oo�o�oGh4Soeo�o8�o<�oEj5�o�'� K�o�