��   u�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����PASSNAME�_T   0 �$+ $~'WORD  ? �LEVEL  �$TI- OUT�T D&F/�� $SETU�PJPROGRA�MJINSTAL�LJY  $�CURR_O�UwSER�NUM��STSTOP_T�PCHG V L�OG_P NT��N�  6 COUNT_DOWN��$ENB_PC�MPWD� $D�V_� IN� s$C� CRE��MA RM9� T9DIAG9(��LVCHK F�ULLM/�YX=T�CNTD��MENU�AUT�O+�FG_DS]P�RLS�U�F��$$CL(   ���!���	��	 V� I�ON( � �:�$DC�S_COD?�|��%�  WF'�_S  *�� $ �&�A91V"!�^ 
 $ !���-�/�/�/�/? ?&?<?J?`?n?�?�?��?�?�?�?�?��#SUP� �+�?O�#�F$O6OvO��  �L�A���O� � �� V�?[t&��j�� �BCO_���G�O�� @ AV6__P