��   L�A��*SYST�EM*��V8.3�382 5/9�/2018 A� 
  ����CELLSET_�T   w�$GI_STYS�EL_P �7T  7I�SO:iRibDiTRA�R��I_INI; ����bU9ART�aRSRPNS1TQ234U5678Q�
TROBQACKSNO�� )�7�E�S��a�o�z2� 3 4 5 6� 7 8awn&GINm'D�&��)% ��)4%��)P%��)fl%SN�{(OU���!7� OPTNA �73�73.:B<;}Ta6.:C<;CK;CaI_DECSNAp�3R�3�TRY1���4��4�PTH�CN�8D�D�INCYC@HG�KD~�TASKOK� {D�{D�7:�E�U: �Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V��Tb@SEGq�T�8�T�@REQ�d��drG�:Mf�GJO?_HFAUL�Xd8�dvgALE� �g�c�g�cvgE� �H�dvgNDBR�H�dg�RGAB�Xtb �F��CLMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVERSION�ix  ��:�$'61�r���p��q�t+ �UP0 �x�Style Se�lect 	  ���q�uReq.� /Echo��N�yAck�����InitiaQt�p�r�s��#��@�O�a�p���	���  ����*������)���������q���O�ption bigt A��p ��B���C���Decis�c�od;��w�pTry�out mL���
�Path s�egJ�ntin.z��8,� cyc:���\�ask O�K!�Manual opt.r�pA"��ΜB"�#�Μ�C"�?�Δdecs�n ِ��pRob�ot inter�lo�"�<� i�sol3�"�̕CҚ�i/�"�x�ment��x�ِ���"���^�statu�s�
	MH ?Fault:��'�{�Aler��ǁ'���p@r 1�z L��[�m�+��; LE_COMN�T ?�y� � ����������ۿ� ���"�4�F�X�j�|� �Ϡϲ���������ƿ@��<�N�`�r��s�25 ��Too�l Change̛ҵ�ap��v�uto C��r{�yߋ��31��Repa�ir2���3&�r�4��Reserved��spY�V�|�� d����������� 0��@�f��߄�Z�� ������������ (O`rH��� ����$J \2l��z�� ���/4/F//W/ |/�/�/v/�/�/�/�/ �/?0?B??߼��? �?�?�?�?�?�?OO ,O>OPObOtO�O�O�O �O�O�O�O__(_:_�L_*�|?ZUZDT� Tes���B�reak��eck R?P?b?�_�_o�_(o &oLo^o4ono�o�o|o �o�o�o �o6H X��x��p���{[(z��E_E�D� ��0��epm�$�Uv	��F�� P��w�a���P�S�����R��������O_Bm�  �����I� ���[� q�J����ӟџ��	��T� ɩ�� � �#�]�o�d������� ��ѯ�����+�=��O� c�a�?� ���LE��  @���/� T_Lɿ���ۿ��,�*�  SS����Rό�� l�������������z\�E�C�i�{����1���1���21����OPmW1ޞ����� �1��E����L_1�#� $��1�$�1���E���~��PTI1ߓߑ������-�~XF.H��\�1��d�$STY�LE_COUNT|�������ޝ�ENAB̀�s������ �� ����'9KU ��k}����� ��1CU_ eq^y���� v���/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f?�x?�?�?�?�? �M�ENU�����6N�AME ?%��(%*DO�}YOSO�>B	PRT03_'R01XO7I$DE�]DS[jC5qO[Om@6�O�Om@7�O�O�O�OiD�9_#_5_G_iC11a_�O�P2�_�_�PpO r_�_5o oYoDo}o�]_�_�Q8�o�o�P`_�ol@20�oouo�o t�_*<���TT  EE��ICG�� ��-�?�Q���u����Q[3�_z~D�VREGPR2��|��3���X���4-�]�ER`BO{�>O����RG��˟  �ʃ�o��̼�P���OB�  ^�jB4Џ\� h2�[� o��4��Я	��p10���O���P�� J���F���.\�]��jB5��`�����!�d�FL�0K��o�m�UPbϛψ^Ͽ�\�p���,��y���� 
!��;�  �*�c�����2ύߦϨ�T�LIM�����'�j�-��LH��$<j�� �� ����v����Z���f�?���G0�i�,���8�1O����~���R�����
��.����"[��J�  ��r����  q����#� 4K�p:s� �fb��q��� �����p-�/� ʈ/;/�p5*/c/� ��R/�/�p@z/�/  #.�/�/�pH�/?� `�/+?��?S?� �B?{?�pX�x�?�'��%�2101_�TC�?��* TCɿ�w�53�?�?�?z~�45@?O)O;O��ZZF7dOvO�O�O7TLD̀N1�@�OJ���F2_�H�"Q#PK RT_��JV+_��I�"T1N#����VK���"rT�_��Q��V�_�YT"T2�_��:fo9LRAo"�뫊fko�"V�o"��"V�o�rV�o��rVQߊ��y�z�  ���VB�328_Z#DT��G�t9��OD��|~B�{�W@�j�D���p���ˏW@⺏ ��p�����
�C��  2�k�W@�Z���V�F����W@�Ȫ��V�xҟ�  A�2�U��"�[��J���V��r����үW@¯�����#�校/J��!�:�s��rb����(���ÿ�a`���0�ڿ����;��7*�c�  q����?zϳ�v�:���Ϟ�����u�l��+ߞ�N��S�v��B�{ߞ�X@jߣ�v���ߝ�_�ߎ��  ���g@
�C��9j��nZ� �������v������
���}��3��)/Z����J����y/���������   �/����I"��?J�i�r��i?�������Ĳ� ������; �*c  ����z�vZ�� ���/v��*/��/S/vIPD/}/��j/�/v�P�/�/��/�/  �P�/?�
?C?09`4?m?� 	�?1!P�?�? 
�?�?0��?O�a@�?3O01�ZOJO�O  rO�O�q@�O�O�@A��O-�OD#_�@�_K_�p5:_s_�@�b_�_�p9��_"�A�_�_�pG�_o�  o;o�pL�*oco&`HRo�o�pQzo�o&`z�o�o~?�o�"d��o+�?O"d� B{O�kD�����o@B���o?��t2�k�>���A������ߏ��ҏ�nO/�
��Z��O~�A�<r���_ϟi��ß���T��"�  g����K� �Po�q�NaE2b��� 1#�_¯����"�Pگ�֠6�;�8���b�  0蟉�"�!x���]R��ۿ_P<