��   Z=�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����SW_ADVFU�NC_T   �P $FAST�FLTREC � $AUTO_�REWELDEN�UMN TRIESVE $^YN Ge�MOTION_L�OCKE�&CwELL1 L8 �HOME_POS�_PReSH�P�OLLEPB_N�OQ�STROK�E�SOPRUN�E�IO1t� 7$DO_JT�e�IMANU�A�PRCA�LT 8CLR�XFR XOP�ENCxRE�P|�ATPNCE ������/? >�NOT�AB�$WDE�NB4$/COM�>W!��7*t$�P�RTI��#�R=Q   �(��&MNT�,�#�(O�UTTO�,�(I�WV+ 4I_LV� >576RTHM�F�\6U7PCMPx|6U7MTWS]�6�:LD�;�0�9� ��:�1k'IMINF�z(�3�=� �1cSP=.B'DX� x(KC�#
 !���ONFIG1�, %YWD_C�TLS ��_�6!EQ�GLCH_�FFe 0_TYP�E�BTD_AFT�ER_CD�@DU_MP_CH�$�0_HID��A�F�A�CYCLc�ADE9FZ 	VWDU��A�VENDO�$�PS�@_DSB_-D��$<UE�A�@�TDFFEXCH�ri �BPREV<ERCOUNXP�N C_O�GWAR~�$CUSTOS�o@T�A�@�WOND�LY�XF�UFRCΝ1NWDH LR�\ CVRS�@I��@SP�AeEXT�_WSD_SCH~UDX_CFG� �PdA$OK2SK�P_SPO�S�QC�NF�FQWKVI�EWd�BSHRTFTnIT�SJ�0IT�SNlPLOaS`T�RNSe�&EQ��� ^T_�GUN�)�d�(ST0tA�j�(|BU�lp"�(Q ~"t�)P|Fs0�(�4`y�(HV�~y�(M�{�q�(@0�)�q��%GO_BINMPV�&�w{y��y�y��"��y�@��{EQ7[��(�`C�P�(��{yD1:����zƂ�]z_BY9P܍�*O�B��i5!^)�OD�ER]G��`PRS��g��(�;����:��/ENW=ɒ76WSOK�'䔻&��F���MW_FLQW��&��C�`Si��H���I��VCL��2���X���똏BUOP��֣˪C�3��G������<:��TCGN�P��`�U�NESA�����H^ �����AIR�3»�HD�h�Ẁ�x��yE7(�76NS�@õ?�?�?�?A�ܚ� ��cSE�TU�p qIY�`TTUDQ�E�VQUDBAC�KU�QVRDROPmO�A%WQPI������2��ӟBCT�RL���#G_SEQUENT��a��Rd� REN��Af'PULC��PTa{`�NT$�OT�PrB�4���a��_�� T_ �UFp�a�@��p��p �_IDX�$SOF6=OUa �����@TISp���q�h��ӫ��P��"�DEcLA�Sb�3�QU�vWOS�WCU�cqO[�qk�MUL�� a���Z��!G����EQ�P��Vt@MBa4g�cb���AF���P�@s AT�EP�B4� G�S��A@�	�EV�/�H	��E �O�D��pC� �|k�"h� x�Fp}�S�o���|� k�X�T �����R��j�Q��` GG:���OO�@G�abS�}�g �p�36�Bg��È�ƦFT��ixGN�hPED��A�C+LS�cM��L�0�u�1�N�@ ��`M�� ;�B���O�I�Q_�PARA%c`�O�C_NAMZ�	y$/P_�4PAU��������uA , ��CO��!LF~  �kA��A�c� �$_MAJOR�@GcL @�EO+�h�Or`$U�A��%SSD�Xր�R1�@o@h�@D0I�ME��M_FA�A>�ST�A2"<�t g =MEDLA���D��_�#0��P$I�f�0LVLV"�ARL��`�c@�_����K+@*T�ARI3TYf�1SO���*[��p`Ea��&[�_�!Pr`3F 4��D�!��@!3�')�OH@4�7Tg��̘`4��#x;[�USGER12G�3�:2�;2V9ART�8�4�;8�8�4w7EFE�#��`C}��҆99FWW#|TL[�MDSON�Ȍ|DsITW�K[�AcLH���D[�OP?K��DW7HX�aH�D=�A!P!.�Sw7Qaх8�=S[�E��AX\T[�I�NRQT+�vZ78IcNI9�S[�WD���O̐ �W��Z5KCH	��Z�&z�(�Tݖ �+fݗ�Pi!4l3h^I�Zf3hB9zfݖ�AL1Mbǜd�gIN�k�c ݖW!�6�e�j�6�e3iP�7vݖA�h8s/z8�hVsݗCFL!hts`k{y�sݖ"�AR�h<�tݖAHDBS�c�D�t�yM i�t�hI i�gOTO�h0��w�AUT�FL��wCROV��l��$�1AU@��S�0@W���gA>P�Q�h̓ÉX�ݖTppЉ�gNRD�W*���vpCO�&J��T�����#$LEA@���Tw��V�qK��x�x��SDEV_N��p�T���йNDXK� �ә�DX�J�3Ca
>��
��WC��p.��T/��ACC��z_�Cc���$���A�� ����o�  � w�d�VE�RSIQm��  �:�$�SPOTADVF�=�  o�#w�����{���CELL ��d��{�ϧj�ܭ���{��D�;�M�CtI�c�Ga� a�A��f�������Fw���a���ܿ� ��Sim info�rm:����Ha�
�=��ϤONFIG ��z�����κ�� ����[EP��7���2�5�π�ρ̾�ʡ|�Ϥ
O�M  ��� �������p߂�Q�EQvj�1ܫȹ� ����������%�7�I�[�m������ ���������
��.� @�R�d�z�r�ߎ�j� |���������"4 FXj|���� ���0��d ��`������� �//,/�� �J/t/ �/�/b/�/�/�/�/? ?����<?n��FL �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�Ov?0_Z?_ V_h_z_�_�_�_�_�_ �_�_�/oo@oRodo .opo�o�o�o�o�oD? F_:_�?�? _r� �������� &�8�J�\�n������� ��_2_D&�o"�4� F�X�j�|�������ğ �oП������<� f�x��������� ���j �>�P�b�t� ��������ο��� �(�:�L�^�pς��� �������� ��$� 6�H�Z�l�~ߐ�R��� �����ߴ����2�D� V�h�z�ܯ����Ϙ� 6���
��.�@�R�d� v��������������� *<N������$SPOTEQ�SETUP 1������ �� %$*����@/S>g
�ȔE,���h���[�z����/#+ ���� L"�~�A�  @] $/�t"e/w/�/+/h�/n���#�|$�/�d4�(3��	�-��	? ���t? ?�?�?�?�?�?�?m ����/��/�O �O�O3/E/W/�/�/_ _�OO_�/�/Og_? /?A?S?e?o�?2oo VoAoSo�oOO+O=O OO�osOU_#5G�O �O�O3_���[� o_�_�_��_�_�_�_ �_��sȍ����ۏ� &��o�o�o�o�o7� ���ϟ�gy�� /�A�S�韏�	��-� ?�Q�c�u�����B�� f�Q���u�������M� _�q���������W�i� {���%�g������� ��)ϣ���ǯٯ������TAT 1�	 ��<$ڙ��� a�����F��j�e�S�}�������NUMEQ  �?�W��WELDIO 1�
�ظ߼Ѫ���c��P�  ���x
}��ћ��� ������	�'���� .@R��n	+���������+�85
0aC
u[�
����� �����uN�d�v��� ��\f/x/�/���/ �/�/�/?rt>?P? b?t?�?�?�?�?&�? �?\�?��SO�wO �O��/"/4/F/ ? _$_6_�/�/l_~_�_ �_�__0?�_�_o o 2oDoVoho�?�o�oO O,O>O�obO#5�O �O�O�O�O�O�_�� �L_^_�*�<�N�`� ��_������̏ޏ�� ��~o(�J��o�o�� �o��>���DVh z����j�|���� 
���֯����^�(� ��T�f�x��������� Z�Կ��`�r�,ϖ�W� i�̟�����&�8� J�4��(�:�L߶�ȯ �ߔߦ߸�"���6� � �$�6�H�Z�l�~�� ���ϸ�B���x� 9�K������������ �������b�t�.@ Rdv���߬�� ��*��N` ��d��0��$��� Z�l�~���������/ �/�/ �/�/�/? "?t/�X?j?|?�?�? �?�?�?@�?Ov� ��mO�bO�O// */</N/`/:?,_>_P_ �/�/f_�_�_�_�_ _ J?oo(o:oLo^opo �oO�o�o"O4O�oXO +�OO�O�O�O�O �O_�_�_���x_ �_D�V�h�z�����o ԏ���
��.�@� �od��o�or�şן :��ޟpx