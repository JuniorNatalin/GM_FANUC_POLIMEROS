��   �=�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����EIP_CFG_�T   � �$VENDOR � $DEVT�YPE>PRDC�ODIREVIS�ION>FAST�_UDP 5 K�EEP_IO_A�nSCNpOPT�` Sp $LOAgDED� �CC� �IG�ED_MO�D�NET�EX�PLCIT_MS��$HIGH_�SPEE�$E�N8021pDS+CP� Hp �� �SPARE���&ONN. |� $HOS� �!B SC9ENA�BL$STA�TN _SZ�S�^TOAPI�OETrIgA�R]�V�BW&Mo��&SC.�  7�CXQ�[XX_���CX_��[ kRs�)%'FLA�MU�L�TR�� C_�O�["TOD&IC$i �AS�Z 'sEC{#�#TIMV�CN� Z�&PAT�  @$IDA_FORMA���!�&� �"9"FIG�^�"2�+�!�$ANALOGI� o  4OU� f8FM�$Q�(� �$$CLA�SS  ����e1��.��.Z0V�ER_c7  �:�$'�0 �8. d��D��0�0> �?�3���7/ ��4(� 2�;@ p!�124.11.�240.31 �xh���� 04���!C�ell ctioCn1�?���1�12_D�<gD�:!l1�O��!?Conne:BbA@�O�OKOyO�O�O3_ 1_C_�Og_
_<@*E�_ �_K_]_�_�K5�_o #o�_Go�_<@6Qo�o �o6o�oZo<@7�o�o �o'�o<@81a s�:<@9�� ����<@A�A� S��w��<@B���� Ïf�珊�<@C�!� 3�֏W���<@Da��� ��F�ǟj�<@Eџ� ���7�ڟ<@FA�q� ��&���J�<@G��� 󯖯���<@H!�Q� c����*�<@I���� ӿv�����<@J�1� C��g�
�<@Kqϡ� ��V���z�<@L��� #���G���<@MQ߁� ��6߷�Z�<@0����0�ߨ�)���nO1�a� s���:�<@P���� ������<@Q�A� S���w��<@R���� ��f�����<@a0#0����Y��nTa� �F�j<@U���192.1�68.1A=�BO�utputVlv	#<QN�8�;�� LW����	U �B��0�g@��PRT38_R0s1 )"g@d!�A3_K/]/ 2�_�?
MH InX^ o}�,�_�-�O/? �/�/6oo�-:/�?B? ��?�4#�oOO / AO�?6!O{O�O0O�O TOfA��O�O�O!_�Of@401_\_n__�_ 5_GP�/�_�_�_o�_ FQ?;oMo�_qooFQ �?�o�o`o�o�oFQ�/ -�oQ�oFQ�/� �@�dFQl?�� �1��FQ�?k�}� � ��D�FQjOۏ폐�� ��FQ�OK�]� ���$��f@5J_��͟p�UN�NINϡ	PE�ND��	ERRO�򄣔�_+�=� ��a�����*o����P� ѯt����o��p/2�5
��DKL C?hangerQ�r +�ɯ����z �����!�Ŀ���[� m�ϑ�4Ϧ�Z����� ��ߤϦ�ʏ;�M��� q�ߦ�:��߽�`�����f@6���-���Q� �������@���d� ኯ�����1���� ��k�}� ���D��L���������$EIP�_SC 2����. @�����.!N����[@]���!}����� ,>Pbt�� �����//(/:/L/^/���:�/t/ �/�/�/@Rdv'? 9?K?�o?��?�?�? �?�?�?�?O#O5OGO YOkO}O�O�O�O�O�O �O�O�/__C_U_g_ y_�/�/?�_�_�_X? �_|?-o?oQocouo�o �o�o�o�o�o�o );M_q��,_ >_������_�_ �_�_m����ooǏ ُ����!�3�E�W� i�{�������ß՟� ����/�A��e�T� ������ �2�D�V�� �+���O�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ����r�����#�5�G� Y�̯ޯ�߳���8� ��\���1�C�U�g� y������������ 	��-�?�Q�c�u�� ߈���������f�x� �ߜ�M_q���ߧ ����%7 I[m���� ���/!/��E/4/ i/{/�/ $6�/ �/?~/?�S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�OR/�O�O__'_ 9_�/�/�/�_�_�_? ~_<?�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CU�O �Ohz���F_X_ j_|_-�?�Q��_�_�� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�� I�[�m�����ǯ ٯ�^����3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛ�2��Ϯ������ ߌ�����a�s߅��� ^����������'� 9�K�]�o����� ���������#�5��� ��H�Z�������&�8� J�\�1�߶�g y������� 	-?Qcu� �����x�/� )/;/M/���������/ �/�/>�/b?%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O/�O�O�O�O�O �Ol/~/�/A_S_e_�/ >_�/�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o�O �O(:o��__ *_<_����_�_G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������X�ԟ 	��-������� �����ϯB���� )�;�M�_�q������� ��˿ݿ���%�7� I�[���nϣϵ��� ��L�^�p�!�3�E߸� �ܯ�ߟ߱������� ����/�A�S�e�w� ������������ ����O�a�s����� 
��������d�v�' 9K]o���� ����#5G Yk}��8��� ��/��������g/ y/�/���/"�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;O�_ONO�O�O�O �O,/>/P/__%_�/ �O�/m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�olO ~O�o�o/AS�O�O �O�O���D_V_� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o������� ɟ۟�`r��G� Y�k�������ůׯ �����1�C�U�g� y���������ӿ��� 	�ϲ�?�.�c�uχ� ����0������x� �Ϝ�M�_�q߃ߕߧ� ����������%�7� I�[�m�����L� ^������!�3��ϸ� ���ύ�����$�6��� ��/ASew ������� +=Oa��t ���@�R�d�v�'/ 9/K/��o/���/�/�/ �/�/�/�/?#?5?G? Y?k?}?�?�?�?�?�? �?�?�OOCOUOgO yO��/�O�O�OX/ �O|/-_?_Q_c_u_�_ �_�_�_�_�_�_oo )o;oMo_oqo�o�o,O >O�o�o�o�O�O �O�Om�__� ����!�3�E�W� i�{�������ÏՏ� ����/�A��oe�T� ������ 2DV� �+��O��s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿr����#�5�G� Y�̟ޟ�ϳ���8� ��\���1�C�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ψ��������fψ���	��4�� $i,�,d��b�t� ���Ϫ��������� (:L^p�� ����� $ ��H7l~��u� '�����/����)/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?U�?�? OO*O�����O �O�O/�O?/�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXo�?|oko�o�o�o��o	�[O�j:�j,hC,gBT�C�o �O������� �!�3�E�W�i�{��� ����ÏՏ����o� �A�S�e�w��ooZI ,ݟ��Ot
�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�����6�ÿ��� ���~���bO��Ɵw� ������ �������� �+�=�O�a�s߅ߗ� �߻���������'� 9�п]�L����� JO<�nO���#�5��� ��k�}����������� ����1CUg y������|� 	�-?Q������ ����B�T��/ )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�? �?�?^p��EOWO iO��O /�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o�?=o,oaoso�o�o 
OO.O�o�o�O �OK]o���� �����#�5�G� Y�k�}�������ŏ\o �؏��1��o�o�o �o������"4ʟ�� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�����r��� ��˿>�P�b�t�%�7� Iϼ�m����ϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� �ߐ���A�S�e�w� ���Ͽ�������h� z�+�=�O�a�s����� ����������' 9K]o���<� �������� ��k}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???�c?R?�? �?�?0BTOO )O�MO�qO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_p?�_�_!o3oEoWo �?�?�?�o�o�o�oHO ZO/ASew �������� �+�=�O�a�s���o ����͏ߏ�dovo�o �oK�]�o��o�o���� ɟ۟����#�5�G� Y�k�}�������ůׯ �������C�2�g� y������"�4���� 	�|�-Ϡ�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ��P�������%�7� ����ο����(� :������!�3�E�W� i�{������������� ��/ASe�� �x���D�V�h� z�+=O����j� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/�#??G? Y?k?���?�? �?\O�1OCOUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_0?�_�_�_�_oo �?�?�?_oqo�o�oO O�o�o�o%7 I[m���� ����!�3�E��_ i�X�������$o6oHo Zo��/��o�oJ�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯v���'�@9�V�f�̇�x�	���4� $�,d,e\�¿ԿG��H�d��'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }���ߐ��������� Ώ���C�U�g�ڿ�� ������������	�� -�?�Q�c�u������� ����������; *_q����,� ������I[ m������ �/!/3/E/W/i/{/ �/�/�/�/Z�/�/? ?/?�����?�? �? 2D�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_�/�_p_�_�_�_�_ N?`?r?#o5oGo�?ko �?�o�o�o�o�o�o�o 1CUgy� �������_� 
�?�Q�c�u��_�_o �oϏ��foxo)�;� M�_�q���������˟ ݟ���%�7�I�[� m������:�ǯ��� �����������i�{� �� ��$�տ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�ԯa�P߅ߗߩ߻� .�@�R���'K� ��o��������� �����#�5�G�Y�k� }�����������n��� ��1CU������ f���F�X�	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/ �/�/bt��I?[? m?���?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _�/A_0_e_w_�_�_ ? ?2?�_�_oz?+o �?Ooaoso�o�o�o�o �o�o�o'9K ]o����N_� ���#�