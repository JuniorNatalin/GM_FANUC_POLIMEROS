��   #L�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETGy �D�HCP_CTRL~.  0 7 �ABLE? $I�PUS�RETR�AT�$SET�HOST�4��DNSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!��* �D $PRIM�AR_IG !$?ALTERN1��<WAIT_TI�A �)��FTޒ @� LOsG_8	�CMO>�$DNLD_F�I:�SUBDI�RCAP�  \q��8 . 4� �H�ADDRT�YP�H NGT1H��	�z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV����PIN�FO.   �$$$XH��RCM+8� ?$| ��QS�IZ�X�� TA�TUSWMAIL�SERV $P�LAN� <$L�IN<$CLU����<$TO�P7$CC�&FR�&��JEC�!�%EN�B � ALAR�!B�TP�/3��V8 S��$VA5R79M ON,6���,6APPL,6PAp� -5B +7POR��#_12ALER�T�&�2URL �}�3ATTAC���0ERR_THRO�3US�9�!�8�R0CH- YDMA�XNS_�1�N1AMOD�2AI� �o 2A� (1APW7D  � LA �0v�ND)ATRYsFDELA�C2@�'`A�ERSI�1A�'R]O�ICLK�HMt0��'� XML+ \3S/GFRM�3T� X3OU�3Z G_��C�OPc1V�3Q�'C8�2-5R_AU�� p� XRN1oUPDX�PCOU�!SFO� 3 
$V�~Wo�@YDUMM�Y1�W2?�RD�M*	T $DI�S���,�SMeB�
"�BCl@bDCI2AI&P�6EXPS�!�P�AR�9��RCL^� <(C�0��SPTM
U� P�WR�h'f �<�Po l5�d�!�"%�7YCC��% 0�fR�0�eP�� _DLV�tf���SNIFF� � �$?�s�_ST�$: G!G�$0q'v�PP��$�@MvBUFF&RPbq��3IF�I��>XPOSAV��dND�!\3� ���0WERUE%�EO+WN��AEa0�dF(e"\�`o3 ��o�bX_`�#Z�_INDE,C%�OZdpE�dUR4�D��F��t�  � t �!�`MO�N�m�D�n�HOU�#EyAt����������LOCA� Y{$N�0H_HE�K�PI"/ 3 $ARP�&�1�vq�W_~ wDEF'�;FA�D�01#��HO_� �R܂EL	% P K Y !�0WOa` -poACCE� LVp�k�2�qK ICE���p ��$*� ? �������%
��
���`S$Q���  ��:�$'0 ј
�
��F����ܐ��w�$� 2�T"����>���� ���!������^���ί��������À_  ���4�F�X�j� |�������Ŀֿ���\��� _FL)p Й��� �����B�����nx�2�����SH)`D 1��d Pᯤ�� ���Ͽ��Ϸ����<� ��H�#�qߖ�Yߺ�}� �ߡ����&�����\� ��C��g����� ����"���F�	�j�-� c������������� ����Af)�M �q�����, �Pt7�[m ����/�:/��3/p/_/�/W/�/��PoPP_L�A1�_x!1.�"0�/�{&�%1?{&25c5.;5�/}#���#2�/
>o0?0?B?T?f63p?
>�0�?�?�?�?f64�?
>_@O O2ODOf65`O
>�@ �O�O�O�Of66�O
>�OP�O_"_4_�RC��G ��������C�� Q�	 �/�^<�_o1oo�UogoyoLo�o�ox(P �o�o�o�o'9K@]����^v�w)�1�1��
Z�DT Statu�se�@�R�d�y'}�iRConnect: irc��//alert� ����ӏ�x�.��%��7�I�[�m�!��P�bb�d��r����� ̟ޟ���&�8�J��\�n����$$c9�62b37a-1�ac0-eb2a�-f1c7-8c�6eb53b4834  (�ӯ&� ��	��-�{%<Qb��X��R^��zP��Plc�
�Q��T,$� ��b��!��ֿ����� �0��T�;�xϊ�q� �ϕ��Ϲ������,��߀ �Q�%�PDM�_�Q	�+�RSMB 
�)�Qd3&���_�����&��_CL�NT 2�� ���R��"��|�U� 4�F��j�|����� �����-��Q�c�B������MTP_CT_RL ��%�� ���tQ���	}���1�U�|��NIFF� �ߺPN�ONEb�  �fr:snif�f.cap�frs:diss���.dg��Ë��t ��v���P�m�Ga��y�����ԁz�6UST�OM m�|̧$�P �$�TTCWPIPg�m��x\�U� TEL�$�%z�Q�{H!T��$/�rj3_t�pde � R!KCL,/�R}�|�E�!CRT�/�y/�/�RZ$!C�ONS�/�
@!s'mon�/Z$