��  Ij�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����SBR_T  � | 	$SVM�TR_ID  $ROBOT9�$GRP_N{UM<AXISQX6K 6NFF3 �_PARAMF	�$�  ,�$MD SPD_L�ITk�&2*o  � �. ��$$CLASS  ���������� VER�SION��  �:�$�'  1 � �T���R-�2000iC/1�25L���  �aiSR22/�4' 80A���
H1 DSP1�-S1��	P0�1.009, � 	� ���΄   ����������������
=��r9�  :!a������ �@H+  �����߻ Y�� � �v# < �����  �����&  �2�&���>A���$j���
"�����&��� �) 	���� ����������ߗ� ��a��G�����{����B� U K� ��� ��5 :?�����'b�
�E/�/�/�/�/����?��3�?C?U?g?��37�X��=�����J���4]��<���\��cxT�p?�?����0B30+/3L2^2fx����������s"�~��%����8 l�� ^���@����� ��*��*����c	�v 5F����;������Y|��+�\, & ����� �8$P|�?������\'�[�Q���r(�c9	�`D 0���o ���#p�"�@��x���Ou_�_�_�_3���_ ?�_�_o��Z���5Y
��@���p����
�8m  ���8u�����p�THoso�4��?0�?�T3^�R"O4OFK�`�bZOlO~G���H=��4�4��K|4�D	 =��,������o(+  , "� �Bu�O������\'��Y^�q��-r(�6_�H_Z_#�5�G�Y��-|h��_����ŏ o������1��o�o VB10J4Q4^�4�o�m:a# ���(����2�`~8	���� 0��� ���w���yF�''nq��`#�5����-�p��� l�8$�E��s����\'����?�	t������5P�!f <�#�S �u�#�>�'  �
�֯ �����	0�D;���fF�k�}��������ſ׿�D�V� j�T5^5������c��Ɵ؟�x��'��������������+ ���\�O`:"�Dn����[X��D	���t
��e+������ʯ�ߥ������-
(��H��� #�5�G�Y�k�}���L��� "�T6^6F�X�j���r�ϔ϶����	���`�����ϡ��� >0 �������
S�M #\'
��a���t	�� r!��h�z���Ugy�3���������"4FX������Z��n�n���	�� ����//&/8/ J/\/n/�/�/�/�/�/@�/�/�/?"?2<�2? V?h?z?�?�?�?�?�? �?�?
OC�~(O� ���O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_@?o o,o>oPoboto�o�o �o�oOJO<O`OrO :L^p���� ��� ��$�6�H� Z�l�~����_��Ə؏ ���� �2�D�V�h� z��o����0�� 
��.�@�R�d�v��� ������Я����� *�<�N���r������� ��̿޿���&�8� ����P�ʟܟ��� �������"�4�F�X� j�|ߎߠ߲������� ���h�0�B�T�f�x� ����������@�r� d�-��Ϛ�b�t����� ����������( :L^p���� ��� $6H Zl~������ 4�F�X� /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?� �?�?�?�?�?�?OO *O<ONO`O��xO� //�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4o�?Xo jo|o�o�o�o�o�o�o �ohO�O�OU�O�O �������� �,�>�P�b�t����� ����Ώ��<o��(� :�L�^�p��������� ʟ&��\n�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vψ� ������,�>��� *�<�N�`�r߄ߖߨ� ����������&�8� J�\︿������� �������"�4����� ��}����ϲ������� ��0BTfx ������� d�>Pbt�� �����N�/
/ ������p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?" �?�?O O2ODOVOhO zO�O�O�O,//�OB/ T/f/._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�?�o �o�o�o�o&8 J\�O�O�O� __ ����"�4�F�X� j�|�������ď֏� ����0��oB�f�x� ��������ҟ���� �v?�2������ ����ί����(� :�L�^�p��������� ʿܿ�J��$�6�H� Z�l�~ϐϢϴ����� T�F���j�|���V�h� zߌߞ߰��������� 
��.�@�R�d�v�� ������������ *�<�N�`�r������ ���(�:�&8 J\n����� ���"4FX ��j������ �//0/B/��g/Z/ �������/�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OOr :OLO^OpO�O�O�O�O �O�O�O _|/n/_�/ �/�/~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�o�o�o0O�o 
.@Rdv� ��_:_,_�P_b_ *�<�N�`�r������� ��̏ޏ����&�8� J�\�n����o����ȟ ڟ����"�4�F�X� j�������� �� ����0�B�T�f�x� ��������ҿ���� �,�>Ϛ�b�tφϘ� �ϼ���������(� ����@ߺ�̯ޯ�߸� ������ ��$�6�H� Z�l�~�������� ����X� �2�D�V�h� z�����������0�b� T�xߊ�Rdv� ������ *<N`r��� ����//&/8/ J/\/n/�/�/���/�/ $6H?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfO� �O�O�O�O�O�O�O_ _,_>_P_�/�/h_�/ �/?�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $�OH Zl~����� ��X_�_|_E��_�_ z�������ԏ��� 
��.�@�R�d�v��� ������П,��� *�<�N�`�r������� ���߯үL�^�p�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώ�ꟲ������� ����0�B�T�f�x� ��毐�
��.���� �,�>�P�b�t��� �����������(� :�L���p��������� ������ $�߲� ��m���ߢ��� �� 2DVh z������� T�
/./@/R/d/v/�/ �/�/�/�/�/>?�/ t��`?r?�?�?�? �?�?�?�?OO&O8O JO\OnO�O�O�O�O/ �O�O�O_"_4_F_X_ j_|_�_�_??�_2? D?V?o0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�O� �������(� :�L��_�_�_���_o ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �|2�V�h� z�������¯ԯ��� 
�f�/�"��������� ������п����� *�<�N�`�rτϖϨ� ������:���&�8� J�\�n߀ߒߤ߶��� D�6���Z�l�~�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt��� �߽�*��( :L^p���� ��� //$/6/H/ ��Z/~/�/�/�/�/�/ �/�/? ?2?�W?J? ����?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O_b/ *_<_N_`_r_�_�_�_ �_�_�_�_l?^?o�? �?�?no�o�o�o�o�o �o�o�o"4FX j|���� _� ���0�B�T�f�x� �����_*oo�@oRo �,�>�P�b�t����� ����Ο�����(� :�L�^�p�������� ʯܯ� ��$�6�H� Z����r�����ؿ ���� �2�D�V�h� zόϞϰ��������� 
��.ߊ�R�d�v߈� �߬߾��������� ����0謹��ο��� ����������&�8� J�\�n����������� ����H�"4FX j|���� �R� D�h�z�BTfx �������/ /,/>/P/b/t/�/�/ ���/�/�/�/??(? :?L?^?p?�?��?�? &8 OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_�/ z_�_�_�_�_�_�_�_ 
oo.o@o�?�?Xo�? �?�?�o�o�o�o *<N`r��� ������p_8� J�\�n���������ȏ ڏ�Hozolo5��o�o j�|�������ğ֟� ����0�B�T�f�x� ���������ү��� �,�>�P�b�t����� ���Ͽ¿<�N�`�(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~�گ�ߴ����� ����� �2�D�V�h� �ֿ���������� 
��.�@�R�d�v��� ������������ *<��`r��� ����p�� ��]������� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ D�/?0?B?T?f?x? �?�?�?�?�?.�?�? dv�PObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_? �_�_�_ oo$o6oHo Zolo~o�oO�?�o"O 4OFO 2DVh z������� 
��.�@�R�d��_�� ������Џ���� *�<��o�o�o���o�o ��̟ޟ���&�8� J�\�n���������ȯ گ����l�"�F�X� j�|�������Ŀֿ� ��V��ό�����x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���*�����(� :�L�^�p����� 4�&���J�\�n�6�H� Z�l�~����������� ���� 2DVh z��߰���� 
.@Rd���� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? �J?n?�?�?�?�?�? �?�?�?O"O~GO:O ����O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_R? o,o>oPoboto�o�o �o�o�o�o\ONO�orO �O�O^p���� ��� ��$�6�H� Z�l�~�������o؏ ���� �2�D�V�h� z����o՟0B 
��.�@�R�d�v��� ������Я����� *�<�N�`���r����� ��̿޿���&�8� JϦ�o�b�ܟ� ��� �������"�4�F�X� j�|ߎߠ߲������� ����z�B�T�f�x� ������������� ��v� ��ϬϾφ��� ����������( :L^p���� ��8� $6H Zl~����B� 4��X�j�2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? ��?�?�?�?�?OO *O<ONO`OrO��O�O //(/�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFo�? jo|o�o�o�o�o�o�o �o0�O�OH�O �O�O������ �,�>�P�b�t����� ����Ώ����`o(� :�L�^�p��������� ʟܟ8j\%��� Z�l�~�������Ưد ���� �2�D�V�h� z��������¿��� 
��.�@�R�d�vψ� �����ϲ�,�>�P�� *�<�N�`�r߄ߖߨ� ����������&�8� J�\�n�ʿ������ �������"�4�F�X� ����p���������� ��0BTfx ������� ,��Pbt�� �����/`��� ��M/�����/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? 4�?O O2ODOVOhO zO�O�O�O�O/�O�O T/f/x/@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�? �o�o�o�o&8 J\n��O�O�_ $_6_��"�4�F�X� j�|�������ď֏� ����0�B�T��ox� ��������ҟ���� �,����u��� ����ί����(� :�L�^�p��������� ʿܿ� �\��6�H� Z�l�~ϐϢϴ����� ��F���|�����h� zߌߞ߰��������� 
��.�@�R�d�v�� ����������� *�<�N�`�r������� $����:�L�^�&8 J\n����� ���"4FX j|������ �//0/B/T/���� ���/��
�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O �:O^OpO�O�O�O�O �O�O�O __n/7_*_ �/�/�/�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�o�o�o�oBO 
.@Rdv� ����L_>_�b_ t_�_N�`�r������� ��̏ޏ����&�8� J�\�n������� ȟ ڟ����"�4�F�X� j�|��
��ů �2� ����0�B�T�f�x� ��������ҿ���� �,�>�PϬ�bφϘ� �ϼ���������(� :ߖ�_�R�̯ޯ�� ������ ��$�6�H� Z�l�~�������� �����j�2�D�V�h� z��������������� t�f��ߜ߮�v� ������ *<N`r��� ��(��//&/8/ J/\/n/�/�/�/ 2 $�/HZ"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO ��O�O�O�O�O�O_�_,_>_P_b_�%�$SBR2 1�%��P T0 �� ��/�'  �_�_�_�_oo&o8o Jo\ono�o�o�o�o�_ �_�o�o"4FX j|������o �o�o�0�B�T�f�x� ��������ҏ���� ���P�b�t����� ����Ο�����(� :��^�A��������� ʯܯ� ��$�6�H� Z�l�O���s���ƿؿ ���� �2�D�V�h� zόϞρ�j_������ ��&�8�J�\�n߀� �ߤ߶����ٸ���
� �.�@�R�d�v��� �������������*� <�N�`�r��������� ������&
�6 \n������ ��"4FX< |������� //0/B/T/f/x/�/ n�/�/�/�/�/?? ,?>?P?b?t?�?�?�? �?�/�?�?OO(O:O LO^OpO�O�O�O�O�O �O�O�?_$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o_DoVohozo �o�o�o�o�o�o�o
 .@R6ov�� �������*� <�N�`�r���h���� ̏ޏ����&�8�J� \�n�����������ڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� �^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�Pߐ��������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� ������* <N`r���� ���/�&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?/X?j? |?�?�?�?�?�?�?�? OO0OBOTO8?J?�O �O�O�O�O�O�O__ ,_>_P_b_t_�_jO�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�_ �o�o $6HZ l~������ �o� �2�D�V�h�z� ������ԏ���
� � �@�R�d�v����� ����П�����*� <�N�2�r��������� ̯ޯ���&�8�J� \�n���d�����ȿڿ ����"�4�F�X�j� |ώϠϲϖ������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� �������������:� L�^�p����������� ���� $6�F l~������ � 2DVhL �������
/ /./@/R/d/v/�/�/ ~�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�/�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O�?"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0o_Tofoxo�o �o�o�o�o�o�o ,>PbFo��� ������(�:� L�^�p�����x��ʏ ܏� ��$�6�H�Z� l�~������������ ��� �2�D�V�h�z� ������¯ԯ�ʟ�� �.�@�R�d�v����� ����п������� <�N�`�rτϖϨϺ� ��������&�8�J� .�n߀ߒߤ߶����� �����"�4�F�X�j� |�`ߠ���������� ��0�B�T�f�x��� ������������ ,>Pbt��� �����(: L^p����� �� //�6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?(/h?z? �?�?�?�?�?�?�?
O O.O@OROdOH?Z?�O �O�O�O�O�O__*_ <_N_`_r_�_�_zO�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�_ �o�o"4FXj |������� �o�0�B�T�f�x��� ������ҏ����� ,��P�b�t������� ��Ο�����(�:� L�^�B���������ʯ ܯ� ��$�6�H�Z� l�~���t���ƿؿ� ��� �2�D�V�h�z� �Ϟϰ��Ϧ�����
� �.�@�R�d�v߈ߚ� �߾����������*� <�N�`�r����� ����������
�J� \�n������������� ����"4F*�V |������� 0BTfx\ ������// ,/>/P/b/t/�/�/�/ ��/�/�/??(?:? L?^?p?�?�?�?�?�? �?�/ OO$O6OHOZO lO~O�O�O�O�O�O�O �O_�?2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@o$_dovo�o�o �o�o�o�o�o* <N`rVo��� �����&�8�J� \�n��������ȏڏ ����"�4�F�X�j� |�������ğ������ ��0�B�T�f�x��� ������ү���ڟ� ,�>�P�b�t������� ��ο����(�� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� >�~ߐߢߴ������� ��� �2�D�V�h�z� ��p߰���������
� �.�@�R�d�v����� ����������* <N`r���� �����&8J \n������ ��/"/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?T?8/x?�? �?�?�?�?�?�?OO ,O>OPObOtOX?j?�O �O�O�O�O__(_:_ L_^_p_�_�_�_�O�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�_ �o 2DVhz �������
� �o.�@�R�d�v����� ����Џ����*� <�N�