��   ��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ������IA_ELEM�_T   D�$USE  �$LINK_NuOD HTYPC�$SHA\IZ�]DATA  �   d/H�AND7 < {$3 2 � �SLDISTD $COMMEN� �$DUMMY�3D �4�� ��$$CLASS ? �������"��"� VERS�ION�  �:�$�� 2�"�� 
  E0��c��4 ~   C��1rUg�@����/��
/ � '�V/9/K/]/ o/�/�/�/�/�/�// #/5/?d?G?Y?k?}? �?�?�?�?�?�??1? OOrOUO�OyO�O�O �O�O_�O&_-O?O_ #__c_�_�_�_�_�_ �_�_�_4o;_M_o1o oqo�o�o�o�o�o�o �oBIo[o-�! ������� �P�Wi;���/��� Ώ��ÏՏ�(��� S�^�w�I���=���ܟ ��џ���6��+�a� s���W��������ͯ ���D�'�9�o���n	NUM V�    
