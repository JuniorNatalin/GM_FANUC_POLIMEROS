��   R��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����MN_MCR_T�ABLE   �� $MACR�O_NAME %$PROG@�EPT_INDE�X  $OP�EN_IDaAS�SIGN_TYP�D  qk$M�ON_NO}PR?EV_SUBy a �$USER_WgORK���_L� �MS�*RTN � &SOP�_T  � {$�EMGO�}�RESET��MOT|�HOL�l��12�SwTAR PDI �I9GAGBGC��TPDS�RE�L�&U� �� �EST��^�SFSP�C����C�C�NB���S)*$8*$3�%)4%)5%)6%)7�%)S�PNSTR�z�"D�  �$$�CLr   �S���!����� VERSION�(�  ��:�:LDUIM�T  ��� �����$MAXDR)I� ��5
�$.�1 �% � d%��]?���K?�?���" �� �s?�?o?�?�?�?O �?>OPO�?O�O5O�O YOkO�O�O__�O�O L_�Op__1_�_�_�_h�_�_�T! F0 POUNCE�_:�R FRP�!:o���q���R�S �%MOVE TO "yo(fm`#�ob��r^a\c�S.c�E I/O�o�Z�!_I�oIlYf �fE�_i�_�_� N�r����/� ��e������J�\� я��������+�ڏ=� a��"���F���j�|� ����'�֟�]�� ��0�B���ɯx���&�� ��/� �T� �edD���@���d�v� 뿚�Ͼ�п
�W�� {�*�<ɅϽ�ܯ�ϐ� �����;�����߃� 2ߧ�V�h��ߌ��� ����I���m��.�� R�������f�3� ��8�A�{�f���N�`� ������������A�� e&�J�n� ��+��a q�FX�|�� �'/�$/]///�/ B/�/f/x/�/�/�/#? �/�/Y??}?,?>?x? �?t?�?�?�?O�?CO �?O>O�O:O�O^OpO �O�O�O_�O�OQ_ _ u_$_6_�_Z_�_�_�_ �_o�_;o�_�_Io�o no�oVoho�o�o�o �o�oI�om.� R�v����3� ��i��y���N�`� Տ��������/�ޏ,� e��&���J���n��� ͟��+�ڟ�a�� ��4�F���ͯ|�񯠯 ��'�֯K����F��� B���f�x�����#� ҿ�Y��}�,�>ϳ� bϰ��ϘϪ����C� ���Qߋ�v߯�^�p� �ߔ�	�����Q����u�$���  T P�OUNCE}�\�T ������	��f�?� �� �u�$���H�Z������������RE�QUEST CO�NTINU����b5 _=I��t!� %SET SEGMEcP
� �_����q�%}5EARLY��T
Et���N�VALID ROqU@ D��NV_i u������� �2/�V///�/�/ M/�/q/�/�/�/?�/ �/?d??�?7?I?�? m?�?�?�?�?*O�?NO �?O�O3O�O�OiO{O �O�O_�O�OJ_\_G_ �_/_A_�_e_�_�_�_ o"o�_Fo�_o|o+o �oOoao�o�o�o�o��oB�ofx'���� ER I-ZOnQ	� RI�p��
��%EXIT ������� x��ߜ����ҏ���� ����>��b��#����G���Ο}���A���ICK���_3PK���rU����DROP ��$�D�Rq�;�T���SER1Vd�v�$�SVկ;����%DIE �AV RMT A�CT4�]vRT_Ah�ԟ�	��AR��۬N�����w
��
������`������T��OPϯ�s�ٶ�CH�� OPRES������Q�e�v<ÊMH� FAULT R�ECOVR,��?FLT_MH����H���G� CYCLE RATί��#��sM%Rec� Path StgartU�UAE��gSTA�߯�4i�>{�Pause�ߝ��PAU�߿�h��%}}�Resum��Н�[�Y��1�%�}�End���EN�D���سRDo� Bwd Exi��߱�	DOBWD��!����^rom�pt Box Y<3�C�OMPT|�e��+~Pr�yw�Ms�g������OϮ�n�F�z�List M�enu4�LIS�T� �%cpt�atus=U~TA�TPAGH߲�,p�.��try�X{P�ERe��cplear User��1gS�]vĠCL��A>S orcej| Ġ���c</_`/ /!/�/E/�/�/{/�/ ?�/&?�/�*��i?����?<?��ECHO OPTI3��{�0 �0�?�ː����?2OO VO�?O�O;O�O_OqO �O�O�O_�O�OR__�v_�_7_1�Gripx�Љ�2�GRIP�0�Έ��fse�_2��`��_�Δ�pa Presen on�Q��AoRoޱ`�Check Noo3�Q��NO���o���o%�~`pare t��`ick:�OKTO��7�
-O�f>Iqrocee���e?LR2PRC��fZ�p nz�Turn� ON Vacu�um�9�VACU�UM�?e[v	�%�	�FF�#�5�F���K�Ⳗ|m�Blo�woff��s�BL�OWr���{��%�Set Cur=r�`Valv�:�SETVALV��fZu��
�5���To�olq�R�_TOO�L��w�\��aLOS�E `� 1՟�xS_VLE	���X�ޱ �����29��m���$�sޱW��3���Dѯ��ٶuS\�4���5���<�!��5Pe������=�"/�OPE��Y~PN(�~�)�j����~x�*K�ίo��~ܷ+��2���U���M�,ߖ�7߹����M�-/1� CAN 1���*�� N��a���!��2��� ]�'�}����/��?�� �_�/���%�I���
������������aL� p�T�����
��pP�� �I0�mT���R������������_OF ��{���a6og����0��Vk�mS�a7�gHMI �=a �o��
p_HDSRP�gYtl�� ��Ex����Po,��"!���2|˃GET C�URR TL TsYPd���TL_� �T�Vk�%CHECK ő�/�-�HK�/u� �>pMA�TC�� 1DATA�5?�']2q?���o�%
L^6�?�,�2�?jV�8].v,v`UN �?8O�"%@�?��" � aO�O��O�j�$0�#?PRESEN=/�''PRS�O����O `_�O�_�O��_i_�_ �_�_�_&o�_Jo�_o �o/o�o�oeowo�o�o �o�oFXC|+ =�a����� �B���x�'���K� ]���䏓����ɏ>� �b�t�#�5���Y�Ο�}������(��M_T���r�!����W� ̯{�����ï8�節\���������ȿ �POS{����ٱR9F�,� $޿��eϱ�Wϐ� LI�NC�U��ϴ�H <���� R_E�Ϲ��.�ٱC_�X� N�T_�ߒߴ�_T9O�߼� E_z�����߳�TI���  �SM���Xﲲ$J<K�� $C7�I�p������ T2��8��!���	$D�L� BA�����3�w��� OM
�t�����RA��7�B���M�<� 
?x UE�n��BROBOT ?BYPASSq��$SV%RM�|���INTsU�b�BT AUTiO�� j0%�N�LLp<S�1c7�$MACRO�0�XNU|������kSOP�ENBL �������22�����PDIMS�` z���S�U��TPDSB�EX  ��
kU��e/��/ �.