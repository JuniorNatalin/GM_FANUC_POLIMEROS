��   R��A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����MN_MCR_T�ABLE   �� $MACR�O_NAME %$PROG@�EPT_INDE�X  $OP�EN_IDaAS�SIGN_TYP�D  qk$M�ON_NO}PR?EV_SUBy a �$USER_WgORK���_L� �MS�*RTN � &SOP�_T  � {$�EMGO�}�RESET��MOT|�HOL�l��12�SwTAR PDI �I9GAGBGC��TPDS�RE�L�&U� �� �EST��^�SFSP�C����C�C�NB���S)*$8*$3�%)4%)5%)6%)7�%)S�PNSTR�z�"D�  �$$�CLr   �S���!����� VERSION�(�  ��:�:LDUIM�T  ��� �����$MAXDR)I� ��5
�$.�1 �% � d%��]?���K?�?���" �� �s?�?o?�?�?�?O �?>OPO�?O�O5O�O YOkO�O�O__�O�O L_�Op__1_�_�_�_h�_�_�T! F0 POUNCE�_:�R FRP�!:o���q���R�S �%MOVE TO "yo(fm`#�ob��s�S^a�S.c�E I/O�o�Zf!_I�o��rYf�fE�_i�_�_ �N�r���� /���e������J� \�я��������+�ڏ =�a��"���F���j� |�����'�֟�]� ���0�B���ɯx��L���� ��/� � T��edD���@���d� v�뿚�Ͼ�п
�W� �{�*�<ɅϽ�ܯ�� �Ϯ����;������ ��2ߧ�V�h��ߌ�� �����I���m��.� ��R�������f� 3���8�A�{�f���N� `�������������A ��e&�J�n ���+��a q�FX�|� ��'/�$/]/// �/B/�/f/x/�/�/�/ #?�/�/Y??}?,?>? x?�?t?�?�?�?O�? CO�?O>O�O:O�O^O pO�O�O�O_�O�OQ_  _u_$_6_�_Z_�_�_ �_�_o�_;o�_�_Io �ono�oVoho�o�o �o�o�oI�om. �R�v���� 3���i��y���N� `�Տ��������/�ޏ ,�e��&���J���n� ��͟��+�ڟ�a� ���4�F���ͯ|�� ����'�֯K����F� ��B���f�x����� #�ҿ�Y��}�,�>� ��bϰ��ϘϪ���� C����Qߋ�v߯�^� p��ߔ�	�����Q����u�$���	AT ?POUNCE}���gAT����q���g��c�<���� E�}�,���P�b�������������%RE�QUEST CONTINU����5 �_=I��u�� �%SET SEGGMEc�� _�l���r�%5�EARLY�T
E�t��%IN�VALID RO!U@ D��a_iu��s�����v�� ��3/�W///�/ �/N/�/r/�/�/�/? �/�/-?e??�?8?J? �?n?�?�?�?�?+O�? OO�?O�O4O�O�OjO |O�O�O_�O�OK_�O ]_�_0_B_�_f_�_�_ �_o#o�_Go�_o}o ,o�oPobo�o�o�o��o�oC�og(��%� ER I-cZOn�� RI�p���
�%EX�IT����� ��x��ߜ����ҏ ��������>��b� �#���G���Ο}�����ICK����g_PK���tU���DROP ��$��DRq�;�
I���S�ERVd�v�$�SV�կ;���%DI�E AV RMT� ACT4�]vRT�_A�ԟ�	��A�R�۬N�����w

�����`�����T��OP�w
��ޱ��CH�� P'RES�����Q��e�vu�%MH� FAULT R�ECOVR,��?FLT_MH������%G� CYCLE RATί診#�s�%R�ec Path �StartU���EN��STA�߯�4س|n߀�Pause��N��PAU�߿����%}�Resum��ߝ�[�Y��1�%�}�End���E�ND������q�uest Menau��o�5 � U `��w
��%Pro�mpt Box yY3���OMPT|����o�b�myw�M�sg����OϮ�n�߆�Li�L%�LIST8�i��	v%%��tus=<���TPAGH߲�ܠ�z�Op.��tryy���OPERe���<öDo B�wd Exit �agSﵔ	DOB�WD�y��h�:qo�rce User ��r\wĠ�c��c </_`//!/�/E/�/ �/{/�/?�/&?�/�*���i?���?<?��E�CHO OPTI@3� ��0�0�?r:l$ ~?/Oz?SO�?���O8O �O�OnO�O�O�O_�O��OO_�OL_�_4_FS	�Grip�Љ���G'RIP������lease�_��`���_�δ�pa Presen on�Q�Ao�nq�n�Chec�k Noo��Q�N�O���o�j\�B�~`p�are t�`ic9k"KTO��c]�s-O�`rHrr�ocee���eLR�2PRC���;�~�z�Turn ON Vacuum�~��VACUUM�?09�0�B�	�FF�#�5�F��gYy>S�|m�Blowoff��s�BLOWr�叺k���pSet Cu{rr�`Valv�~�ETVALV��fZxHPS5���To�olq�R�_TOO�L��w����`LO7SE `� 1՟�xS_VLE	���mSޱ����29��m�H��>SޱW��3����ѯ�˄�ޱuS\�4@��5����ޱ!��5e������B�|��"��)��N(�~��ܱ)�j����~dcܱ*K�ίo��~,sܱ+��2���U�~�cܱ,ߖ�7�T��~M�-��1�? CAN 1����d1�_ON ϭ�ܷ��<r��2���ϭ�M�������?�_�/���=���������)�_r�ﮋ� LӠrI����wﮋx� �Ө�I0�mT��� R�����������������kX�ܱ6�og����0�kzM�7�gHMI =a� �o��
p_HDR�P�gYu �<PڏT6`���P�o,X�"!�����˃GET CU�RR TL TY�Pd���TL_� T��v��o>pCHECcK ő�/�-HK�/�gY�xdo>pMA�TC�� 1DATA3?�na�"]2n?jV�TIMxI?%
1L^6�?y5  �"�2|�?jV
  x�?�%UN�?�=EM�"%@�?hXSTExp���k^O�OT"/�O�O OT"�q�$0~�#PRESEN=/�  	 �"PR	S�O[xV�zM�D&_��� jpW_��ER�IFYT_\xQVRFY�_�_�_o+o� Oo�_o�o<7�{o�o couo�o5o�o�oD�Vz);��w ���q�p����q��D���z�dt6�y�o��� U@[� m��e��Ǐ<��].S7�p��1����� ��ԟ V�ER�����B1$���8��1���r���ALIc��� � O�a��֯��_ACǯ � �$F��ů:���R8��b��� 	�)�Ğ�}1��ǿ��HI{����A2 �,�P!$߿�f�G�Wϐχ REN�T�����LAY���ϵP����-�F�LT�X��ߘߒ�M�OR�߼� am����s�$W�߂ � h0����Z���M9D����  y�G��T2�����ߩ���I�_N�L�  �B������$JOw���#�c�u������GRP�� DE�L����N��BRK<?x ASE+�A�ROBOT BY�PASSq�� �%RM����I�NsUb�BT� AUTO�� �LEA%�ۯR�Al�c7�$�MACRO�0XN�U_�����kSOPEN?BL X����l�0	����PD�IMS` z�̦�SU��TPDSBEX�>5�kU��e/� �/�.