��   e�A��*SYST�EM*��V8.3�382 5/9�/2018 A�   ����CELL_GRP�_T   � �$'FRAME� $MOU�NT_LOCCC�F_METHOD�  $CPY�_SRC_IDX�_PLATFRM�_OFSCtDI�M_ $BASE{ FSETC���AUX_ORDER   ��XYZ_MAP ��� �LE�NGTH�TTC?H_GP_M~ a �AUTORAIL�_k��$$CL�ASS  �S����D��DVERSION�  ��:�8LOOR �G��DD8�?���m��Mn,  1 <DY�H8G}~}��D'�82 �����i?/Q/c/5/�/�/�-_ �/�/�/��+�$MNU>A�2"�d  8�i�7����b��4�ݿ5	9nQ?B0�=1D��\D8��D�8�ke?� a?�?�?�?�?�?�?�? OO%OOO9O[O�OoO �O�O�O�O�O�O�O'_ _#_]_G_Y_{_}_�_ �_�_�_�_o�_oGo 1oSo}ogo�o�o�o�o �o�o�o	U?~7NUM  ���>a �p�uTO�OL?#;��fq� � í����
�=C-�\Mv���<ʓ�C�м���?��R�ۖ:�t�c<����KC�IZCz��B��1Mu�;�.�fteqC�i}�H3�3Cy��B���Mo��K������ ɏ�ݏ��)��5�_��C��ATc�C*v�S�e���Q� ��՟�������A�@+�M�w�a����B����~ffB��� ����ﯡ���%��1� [�E�g���{���ǿ��@����ϭ�v�s[�y�00